`default_nettype none
`timescale 1 ns / 1 ps

(* rom_style = "distributed" *)
module lut_logsin(
    input  wire  [7:0] idx,
    output reg  [11:0] value
);

    always @* case (idx)
        8'h00: value = 12'h859;
        8'h01: value = 12'h6c3;
        8'h02: value = 12'h607;
        8'h03: value = 12'h58b;
        8'h04: value = 12'h52e;
        8'h05: value = 12'h4e4;
        8'h06: value = 12'h4a6;
        8'h07: value = 12'h471;
        8'h08: value = 12'h443;
        8'h09: value = 12'h41a;
        8'h0A: value = 12'h3f5;
        8'h0B: value = 12'h3d3;
        8'h0C: value = 12'h3b5;
        8'h0D: value = 12'h398;
        8'h0E: value = 12'h37e;
        8'h0F: value = 12'h365;
        8'h10: value = 12'h34e;
        8'h11: value = 12'h339;
        8'h12: value = 12'h324;
        8'h13: value = 12'h311;
        8'h14: value = 12'h2ff;
        8'h15: value = 12'h2ed;
        8'h16: value = 12'h2dc;
        8'h17: value = 12'h2cd;
        8'h18: value = 12'h2bd;
        8'h19: value = 12'h2af;
        8'h1A: value = 12'h2a0;
        8'h1B: value = 12'h293;
        8'h1C: value = 12'h286;
        8'h1D: value = 12'h279;
        8'h1E: value = 12'h26d;
        8'h1F: value = 12'h261;
        8'h20: value = 12'h256;
        8'h21: value = 12'h24b;
        8'h22: value = 12'h240;
        8'h23: value = 12'h236;
        8'h24: value = 12'h22c;
        8'h25: value = 12'h222;
        8'h26: value = 12'h218;
        8'h27: value = 12'h20f;
        8'h28: value = 12'h206;
        8'h29: value = 12'h1fd;
        8'h2A: value = 12'h1f5;
        8'h2B: value = 12'h1ec;
        8'h2C: value = 12'h1e4;
        8'h2D: value = 12'h1dc;
        8'h2E: value = 12'h1d4;
        8'h2F: value = 12'h1cd;
        8'h30: value = 12'h1c5;
        8'h31: value = 12'h1be;
        8'h32: value = 12'h1b7;
        8'h33: value = 12'h1b0;
        8'h34: value = 12'h1a9;
        8'h35: value = 12'h1a2;
        8'h36: value = 12'h19b;
        8'h37: value = 12'h195;
        8'h38: value = 12'h18f;
        8'h39: value = 12'h188;
        8'h3A: value = 12'h182;
        8'h3B: value = 12'h17c;
        8'h3C: value = 12'h177;
        8'h3D: value = 12'h171;
        8'h3E: value = 12'h16b;
        8'h3F: value = 12'h166;
        8'h40: value = 12'h160;
        8'h41: value = 12'h15b;
        8'h42: value = 12'h155;
        8'h43: value = 12'h150;
        8'h44: value = 12'h14b;
        8'h45: value = 12'h146;
        8'h46: value = 12'h141;
        8'h47: value = 12'h13c;
        8'h48: value = 12'h137;
        8'h49: value = 12'h133;
        8'h4A: value = 12'h12e;
        8'h4B: value = 12'h129;
        8'h4C: value = 12'h125;
        8'h4D: value = 12'h121;
        8'h4E: value = 12'h11c;
        8'h4F: value = 12'h118;
        8'h50: value = 12'h114;
        8'h51: value = 12'h10f;
        8'h52: value = 12'h10b;
        8'h53: value = 12'h107;
        8'h54: value = 12'h103;
        8'h55: value = 12'h0ff;
        8'h56: value = 12'h0fb;
        8'h57: value = 12'h0f8;
        8'h58: value = 12'h0f4;
        8'h59: value = 12'h0f0;
        8'h5A: value = 12'h0ec;
        8'h5B: value = 12'h0e9;
        8'h5C: value = 12'h0e5;
        8'h5D: value = 12'h0e2;
        8'h5E: value = 12'h0de;
        8'h5F: value = 12'h0db;
        8'h60: value = 12'h0d7;
        8'h61: value = 12'h0d4;
        8'h62: value = 12'h0d1;
        8'h63: value = 12'h0cd;
        8'h64: value = 12'h0ca;
        8'h65: value = 12'h0c7;
        8'h66: value = 12'h0c4;
        8'h67: value = 12'h0c1;
        8'h68: value = 12'h0be;
        8'h69: value = 12'h0bb;
        8'h6A: value = 12'h0b8;
        8'h6B: value = 12'h0b5;
        8'h6C: value = 12'h0b2;
        8'h6D: value = 12'h0af;
        8'h6E: value = 12'h0ac;
        8'h6F: value = 12'h0a9;
        8'h70: value = 12'h0a7;
        8'h71: value = 12'h0a4;
        8'h72: value = 12'h0a1;
        8'h73: value = 12'h09f;
        8'h74: value = 12'h09c;
        8'h75: value = 12'h099;
        8'h76: value = 12'h097;
        8'h77: value = 12'h094;
        8'h78: value = 12'h092;
        8'h79: value = 12'h08f;
        8'h7A: value = 12'h08d;
        8'h7B: value = 12'h08a;
        8'h7C: value = 12'h088;
        8'h7D: value = 12'h086;
        8'h7E: value = 12'h083;
        8'h7F: value = 12'h081;
        8'h80: value = 12'h07f;
        8'h81: value = 12'h07d;
        8'h82: value = 12'h07a;
        8'h83: value = 12'h078;
        8'h84: value = 12'h076;
        8'h85: value = 12'h074;
        8'h86: value = 12'h072;
        8'h87: value = 12'h070;
        8'h88: value = 12'h06e;
        8'h89: value = 12'h06c;
        8'h8A: value = 12'h06a;
        8'h8B: value = 12'h068;
        8'h8C: value = 12'h066;
        8'h8D: value = 12'h064;
        8'h8E: value = 12'h062;
        8'h8F: value = 12'h060;
        8'h90: value = 12'h05e;
        8'h91: value = 12'h05c;
        8'h92: value = 12'h05b;
        8'h93: value = 12'h059;
        8'h94: value = 12'h057;
        8'h95: value = 12'h055;
        8'h96: value = 12'h053;
        8'h97: value = 12'h052;
        8'h98: value = 12'h050;
        8'h99: value = 12'h04e;
        8'h9A: value = 12'h04d;
        8'h9B: value = 12'h04b;
        8'h9C: value = 12'h04a;
        8'h9D: value = 12'h048;
        8'h9E: value = 12'h046;
        8'h9F: value = 12'h045;
        8'hA0: value = 12'h043;
        8'hA1: value = 12'h042;
        8'hA2: value = 12'h040;
        8'hA3: value = 12'h03f;
        8'hA4: value = 12'h03e;
        8'hA5: value = 12'h03c;
        8'hA6: value = 12'h03b;
        8'hA7: value = 12'h039;
        8'hA8: value = 12'h038;
        8'hA9: value = 12'h037;
        8'hAA: value = 12'h035;
        8'hAB: value = 12'h034;
        8'hAC: value = 12'h033;
        8'hAD: value = 12'h031;
        8'hAE: value = 12'h030;
        8'hAF: value = 12'h02f;
        8'hB0: value = 12'h02e;
        8'hB1: value = 12'h02d;
        8'hB2: value = 12'h02b;
        8'hB3: value = 12'h02a;
        8'hB4: value = 12'h029;
        8'hB5: value = 12'h028;
        8'hB6: value = 12'h027;
        8'hB7: value = 12'h026;
        8'hB8: value = 12'h025;
        8'hB9: value = 12'h024;
        8'hBA: value = 12'h023;
        8'hBB: value = 12'h022;
        8'hBC: value = 12'h021;
        8'hBD: value = 12'h020;
        8'hBE: value = 12'h01f;
        8'hBF: value = 12'h01e;
        8'hC0: value = 12'h01d;
        8'hC1: value = 12'h01c;
        8'hC2: value = 12'h01b;
        8'hC3: value = 12'h01a;
        8'hC4: value = 12'h019;
        8'hC5: value = 12'h018;
        8'hC6: value = 12'h017;
        8'hC7: value = 12'h017;
        8'hC8: value = 12'h016;
        8'hC9: value = 12'h015;
        8'hCA: value = 12'h014;
        8'hCB: value = 12'h014;
        8'hCC: value = 12'h013;
        8'hCD: value = 12'h012;
        8'hCE: value = 12'h011;
        8'hCF: value = 12'h011;
        8'hD0: value = 12'h010;
        8'hD1: value = 12'h00f;
        8'hD2: value = 12'h00f;
        8'hD3: value = 12'h00e;
        8'hD4: value = 12'h00d;
        8'hD5: value = 12'h00d;
        8'hD6: value = 12'h00c;
        8'hD7: value = 12'h00c;
        8'hD8: value = 12'h00b;
        8'hD9: value = 12'h00a;
        8'hDA: value = 12'h00a;
        8'hDB: value = 12'h009;
        8'hDC: value = 12'h009;
        8'hDD: value = 12'h008;
        8'hDE: value = 12'h008;
        8'hDF: value = 12'h007;
        8'hE0: value = 12'h007;
        8'hE1: value = 12'h007;
        8'hE2: value = 12'h006;
        8'hE3: value = 12'h006;
        8'hE4: value = 12'h005;
        8'hE5: value = 12'h005;
        8'hE6: value = 12'h005;
        8'hE7: value = 12'h004;
        8'hE8: value = 12'h004;
        8'hE9: value = 12'h004;
        8'hEA: value = 12'h003;
        8'hEB: value = 12'h003;
        8'hEC: value = 12'h003;
        8'hED: value = 12'h002;
        8'hEE: value = 12'h002;
        8'hEF: value = 12'h002;
        8'hF0: value = 12'h002;
        8'hF1: value = 12'h001;
        8'hF2: value = 12'h001;
        8'hF3: value = 12'h001;
        8'hF4: value = 12'h001;
        8'hF5: value = 12'h001;
        8'hF6: value = 12'h001;
        8'hF7: value = 12'h001;
        8'hF8: value = 12'h000;
        8'hF9: value = 12'h000;
        8'hFA: value = 12'h000;
        8'hFB: value = 12'h000;
        8'hFC: value = 12'h000;
        8'hFD: value = 12'h000;
        8'hFE: value = 12'h000;
        8'hFF: value = 12'h000;
        default: value = 12'h0;
    endcase

endmodule
