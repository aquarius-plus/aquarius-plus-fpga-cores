`default_nettype none
`timescale 1 ns / 1 ps

(* rom_style = "distributed" *)
module lut_exp(
    input  wire        clk,
    input  wire  [7:0] idx,
    output reg   [9:0] value
);

    always @(posedge clk) case (idx)
        8'h00: value <= 10'd0;
        8'h01: value <= 10'd3;
        8'h02: value <= 10'd6;
        8'h03: value <= 10'd8;
        8'h04: value <= 10'd11;
        8'h05: value <= 10'd14;
        8'h06: value <= 10'd17;
        8'h07: value <= 10'd20;
        8'h08: value <= 10'd22;
        8'h09: value <= 10'd25;
        8'h0A: value <= 10'd28;
        8'h0B: value <= 10'd31;
        8'h0C: value <= 10'd34;
        8'h0D: value <= 10'd37;
        8'h0E: value <= 10'd40;
        8'h0F: value <= 10'd42;
        8'h10: value <= 10'd45;
        8'h11: value <= 10'd48;
        8'h12: value <= 10'd51;
        8'h13: value <= 10'd54;
        8'h14: value <= 10'd57;
        8'h15: value <= 10'd60;
        8'h16: value <= 10'd63;
        8'h17: value <= 10'd66;
        8'h18: value <= 10'd69;
        8'h19: value <= 10'd72;
        8'h1A: value <= 10'd75;
        8'h1B: value <= 10'd78;
        8'h1C: value <= 10'd81;
        8'h1D: value <= 10'd84;
        8'h1E: value <= 10'd87;
        8'h1F: value <= 10'd90;
        8'h20: value <= 10'd93;
        8'h21: value <= 10'd96;
        8'h22: value <= 10'd99;
        8'h23: value <= 10'd102;
        8'h24: value <= 10'd105;
        8'h25: value <= 10'd108;
        8'h26: value <= 10'd111;
        8'h27: value <= 10'd114;
        8'h28: value <= 10'd117;
        8'h29: value <= 10'd120;
        8'h2A: value <= 10'd123;
        8'h2B: value <= 10'd126;
        8'h2C: value <= 10'd130;
        8'h2D: value <= 10'd133;
        8'h2E: value <= 10'd136;
        8'h2F: value <= 10'd139;
        8'h30: value <= 10'd142;
        8'h31: value <= 10'd145;
        8'h32: value <= 10'd148;
        8'h33: value <= 10'd152;
        8'h34: value <= 10'd155;
        8'h35: value <= 10'd158;
        8'h36: value <= 10'd161;
        8'h37: value <= 10'd164;
        8'h38: value <= 10'd168;
        8'h39: value <= 10'd171;
        8'h3A: value <= 10'd174;
        8'h3B: value <= 10'd177;
        8'h3C: value <= 10'd181;
        8'h3D: value <= 10'd184;
        8'h3E: value <= 10'd187;
        8'h3F: value <= 10'd190;
        8'h40: value <= 10'd194;
        8'h41: value <= 10'd197;
        8'h42: value <= 10'd200;
        8'h43: value <= 10'd204;
        8'h44: value <= 10'd207;
        8'h45: value <= 10'd210;
        8'h46: value <= 10'd214;
        8'h47: value <= 10'd217;
        8'h48: value <= 10'd220;
        8'h49: value <= 10'd224;
        8'h4A: value <= 10'd227;
        8'h4B: value <= 10'd231;
        8'h4C: value <= 10'd234;
        8'h4D: value <= 10'd237;
        8'h4E: value <= 10'd241;
        8'h4F: value <= 10'd244;
        8'h50: value <= 10'd248;
        8'h51: value <= 10'd251;
        8'h52: value <= 10'd255;
        8'h53: value <= 10'd258;
        8'h54: value <= 10'd262;
        8'h55: value <= 10'd265;
        8'h56: value <= 10'd268;
        8'h57: value <= 10'd272;
        8'h58: value <= 10'd276;
        8'h59: value <= 10'd279;
        8'h5A: value <= 10'd283;
        8'h5B: value <= 10'd286;
        8'h5C: value <= 10'd290;
        8'h5D: value <= 10'd293;
        8'h5E: value <= 10'd297;
        8'h5F: value <= 10'd300;
        8'h60: value <= 10'd304;
        8'h61: value <= 10'd308;
        8'h62: value <= 10'd311;
        8'h63: value <= 10'd315;
        8'h64: value <= 10'd318;
        8'h65: value <= 10'd322;
        8'h66: value <= 10'd326;
        8'h67: value <= 10'd329;
        8'h68: value <= 10'd333;
        8'h69: value <= 10'd337;
        8'h6A: value <= 10'd340;
        8'h6B: value <= 10'd344;
        8'h6C: value <= 10'd348;
        8'h6D: value <= 10'd352;
        8'h6E: value <= 10'd355;
        8'h6F: value <= 10'd359;
        8'h70: value <= 10'd363;
        8'h71: value <= 10'd367;
        8'h72: value <= 10'd370;
        8'h73: value <= 10'd374;
        8'h74: value <= 10'd378;
        8'h75: value <= 10'd382;
        8'h76: value <= 10'd385;
        8'h77: value <= 10'd389;
        8'h78: value <= 10'd393;
        8'h79: value <= 10'd397;
        8'h7A: value <= 10'd401;
        8'h7B: value <= 10'd405;
        8'h7C: value <= 10'd409;
        8'h7D: value <= 10'd412;
        8'h7E: value <= 10'd416;
        8'h7F: value <= 10'd420;
        8'h80: value <= 10'd424;
        8'h81: value <= 10'd428;
        8'h82: value <= 10'd432;
        8'h83: value <= 10'd436;
        8'h84: value <= 10'd440;
        8'h85: value <= 10'd444;
        8'h86: value <= 10'd448;
        8'h87: value <= 10'd452;
        8'h88: value <= 10'd456;
        8'h89: value <= 10'd460;
        8'h8A: value <= 10'd464;
        8'h8B: value <= 10'd468;
        8'h8C: value <= 10'd472;
        8'h8D: value <= 10'd476;
        8'h8E: value <= 10'd480;
        8'h8F: value <= 10'd484;
        8'h90: value <= 10'd488;
        8'h91: value <= 10'd492;
        8'h92: value <= 10'd496;
        8'h93: value <= 10'd501;
        8'h94: value <= 10'd505;
        8'h95: value <= 10'd509;
        8'h96: value <= 10'd513;
        8'h97: value <= 10'd517;
        8'h98: value <= 10'd521;
        8'h99: value <= 10'd526;
        8'h9A: value <= 10'd530;
        8'h9B: value <= 10'd534;
        8'h9C: value <= 10'd538;
        8'h9D: value <= 10'd542;
        8'h9E: value <= 10'd547;
        8'h9F: value <= 10'd551;
        8'hA0: value <= 10'd555;
        8'hA1: value <= 10'd560;
        8'hA2: value <= 10'd564;
        8'hA3: value <= 10'd568;
        8'hA4: value <= 10'd572;
        8'hA5: value <= 10'd577;
        8'hA6: value <= 10'd581;
        8'hA7: value <= 10'd585;
        8'hA8: value <= 10'd590;
        8'hA9: value <= 10'd594;
        8'hAA: value <= 10'd599;
        8'hAB: value <= 10'd603;
        8'hAC: value <= 10'd607;
        8'hAD: value <= 10'd612;
        8'hAE: value <= 10'd616;
        8'hAF: value <= 10'd621;
        8'hB0: value <= 10'd625;
        8'hB1: value <= 10'd630;
        8'hB2: value <= 10'd634;
        8'hB3: value <= 10'd639;
        8'hB4: value <= 10'd643;
        8'hB5: value <= 10'd648;
        8'hB6: value <= 10'd652;
        8'hB7: value <= 10'd657;
        8'hB8: value <= 10'd661;
        8'hB9: value <= 10'd666;
        8'hBA: value <= 10'd670;
        8'hBB: value <= 10'd675;
        8'hBC: value <= 10'd680;
        8'hBD: value <= 10'd684;
        8'hBE: value <= 10'd689;
        8'hBF: value <= 10'd693;
        8'hC0: value <= 10'd698;
        8'hC1: value <= 10'd703;
        8'hC2: value <= 10'd708;
        8'hC3: value <= 10'd712;
        8'hC4: value <= 10'd717;
        8'hC5: value <= 10'd722;
        8'hC6: value <= 10'd726;
        8'hC7: value <= 10'd731;
        8'hC8: value <= 10'd736;
        8'hC9: value <= 10'd741;
        8'hCA: value <= 10'd745;
        8'hCB: value <= 10'd750;
        8'hCC: value <= 10'd755;
        8'hCD: value <= 10'd760;
        8'hCE: value <= 10'd765;
        8'hCF: value <= 10'd770;
        8'hD0: value <= 10'd774;
        8'hD1: value <= 10'd779;
        8'hD2: value <= 10'd784;
        8'hD3: value <= 10'd789;
        8'hD4: value <= 10'd794;
        8'hD5: value <= 10'd799;
        8'hD6: value <= 10'd804;
        8'hD7: value <= 10'd809;
        8'hD8: value <= 10'd814;
        8'hD9: value <= 10'd819;
        8'hDA: value <= 10'd824;
        8'hDB: value <= 10'd829;
        8'hDC: value <= 10'd834;
        8'hDD: value <= 10'd839;
        8'hDE: value <= 10'd844;
        8'hDF: value <= 10'd849;
        8'hE0: value <= 10'd854;
        8'hE1: value <= 10'd859;
        8'hE2: value <= 10'd864;
        8'hE3: value <= 10'd869;
        8'hE4: value <= 10'd874;
        8'hE5: value <= 10'd880;
        8'hE6: value <= 10'd885;
        8'hE7: value <= 10'd890;
        8'hE8: value <= 10'd895;
        8'hE9: value <= 10'd900;
        8'hEA: value <= 10'd906;
        8'hEB: value <= 10'd911;
        8'hEC: value <= 10'd916;
        8'hED: value <= 10'd921;
        8'hEE: value <= 10'd927;
        8'hEF: value <= 10'd932;
        8'hF0: value <= 10'd937;
        8'hF1: value <= 10'd942;
        8'hF2: value <= 10'd948;
        8'hF3: value <= 10'd953;
        8'hF4: value <= 10'd959;
        8'hF5: value <= 10'd964;
        8'hF6: value <= 10'd969;
        8'hF7: value <= 10'd975;
        8'hF8: value <= 10'd980;
        8'hF9: value <= 10'd986;
        8'hFA: value <= 10'd991;
        8'hFB: value <= 10'd996;
        8'hFC: value <= 10'd1002;
        8'hFD: value <= 10'd1007;
        8'hFE: value <= 10'd1013;
        8'hFF: value <= 10'd1018;
        default: value <= 10'd0;
    endcase

endmodule
