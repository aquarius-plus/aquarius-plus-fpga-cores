`default_nettype none
`timescale 1 ns / 1 ps

(* rom_style = "distributed" *)
module lut_logsin(
    input  wire        clk,
    input  wire  [7:0] addr,
    output reg  [11:0] rddata
);

    always @(posedge clk) case (addr)
        8'h00: rddata <= 12'd2137;
        8'h01: rddata <= 12'd1731;
        8'h02: rddata <= 12'd1543;
        8'h03: rddata <= 12'd1419;
        8'h04: rddata <= 12'd1326;
        8'h05: rddata <= 12'd1252;
        8'h06: rddata <= 12'd1190;
        8'h07: rddata <= 12'd1137;
        8'h08: rddata <= 12'd1091;
        8'h09: rddata <= 12'd1050;
        8'h0A: rddata <= 12'd1013;
        8'h0B: rddata <= 12'd979;
        8'h0C: rddata <= 12'd949;
        8'h0D: rddata <= 12'd920;
        8'h0E: rddata <= 12'd894;
        8'h0F: rddata <= 12'd869;
        8'h10: rddata <= 12'd846;
        8'h11: rddata <= 12'd825;
        8'h12: rddata <= 12'd804;
        8'h13: rddata <= 12'd785;
        8'h14: rddata <= 12'd767;
        8'h15: rddata <= 12'd749;
        8'h16: rddata <= 12'd732;
        8'h17: rddata <= 12'd717;
        8'h18: rddata <= 12'd701;
        8'h19: rddata <= 12'd687;
        8'h1A: rddata <= 12'd672;
        8'h1B: rddata <= 12'd659;
        8'h1C: rddata <= 12'd646;
        8'h1D: rddata <= 12'd633;
        8'h1E: rddata <= 12'd621;
        8'h1F: rddata <= 12'd609;
        8'h20: rddata <= 12'd598;
        8'h21: rddata <= 12'd587;
        8'h22: rddata <= 12'd576;
        8'h23: rddata <= 12'd566;
        8'h24: rddata <= 12'd556;
        8'h25: rddata <= 12'd546;
        8'h26: rddata <= 12'd536;
        8'h27: rddata <= 12'd527;
        8'h28: rddata <= 12'd518;
        8'h29: rddata <= 12'd509;
        8'h2A: rddata <= 12'd501;
        8'h2B: rddata <= 12'd492;
        8'h2C: rddata <= 12'd484;
        8'h2D: rddata <= 12'd476;
        8'h2E: rddata <= 12'd468;
        8'h2F: rddata <= 12'd461;
        8'h30: rddata <= 12'd453;
        8'h31: rddata <= 12'd446;
        8'h32: rddata <= 12'd439;
        8'h33: rddata <= 12'd432;
        8'h34: rddata <= 12'd425;
        8'h35: rddata <= 12'd418;
        8'h36: rddata <= 12'd411;
        8'h37: rddata <= 12'd405;
        8'h38: rddata <= 12'd399;
        8'h39: rddata <= 12'd392;
        8'h3A: rddata <= 12'd386;
        8'h3B: rddata <= 12'd380;
        8'h3C: rddata <= 12'd375;
        8'h3D: rddata <= 12'd369;
        8'h3E: rddata <= 12'd363;
        8'h3F: rddata <= 12'd358;
        8'h40: rddata <= 12'd352;
        8'h41: rddata <= 12'd347;
        8'h42: rddata <= 12'd341;
        8'h43: rddata <= 12'd336;
        8'h44: rddata <= 12'd331;
        8'h45: rddata <= 12'd326;
        8'h46: rddata <= 12'd321;
        8'h47: rddata <= 12'd316;
        8'h48: rddata <= 12'd311;
        8'h49: rddata <= 12'd307;
        8'h4A: rddata <= 12'd302;
        8'h4B: rddata <= 12'd297;
        8'h4C: rddata <= 12'd293;
        8'h4D: rddata <= 12'd289;
        8'h4E: rddata <= 12'd284;
        8'h4F: rddata <= 12'd280;
        8'h50: rddata <= 12'd276;
        8'h51: rddata <= 12'd271;
        8'h52: rddata <= 12'd267;
        8'h53: rddata <= 12'd263;
        8'h54: rddata <= 12'd259;
        8'h55: rddata <= 12'd255;
        8'h56: rddata <= 12'd251;
        8'h57: rddata <= 12'd248;
        8'h58: rddata <= 12'd244;
        8'h59: rddata <= 12'd240;
        8'h5A: rddata <= 12'd236;
        8'h5B: rddata <= 12'd233;
        8'h5C: rddata <= 12'd229;
        8'h5D: rddata <= 12'd226;
        8'h5E: rddata <= 12'd222;
        8'h5F: rddata <= 12'd219;
        8'h60: rddata <= 12'd215;
        8'h61: rddata <= 12'd212;
        8'h62: rddata <= 12'd209;
        8'h63: rddata <= 12'd205;
        8'h64: rddata <= 12'd202;
        8'h65: rddata <= 12'd199;
        8'h66: rddata <= 12'd196;
        8'h67: rddata <= 12'd193;
        8'h68: rddata <= 12'd190;
        8'h69: rddata <= 12'd187;
        8'h6A: rddata <= 12'd184;
        8'h6B: rddata <= 12'd181;
        8'h6C: rddata <= 12'd178;
        8'h6D: rddata <= 12'd175;
        8'h6E: rddata <= 12'd172;
        8'h6F: rddata <= 12'd169;
        8'h70: rddata <= 12'd167;
        8'h71: rddata <= 12'd164;
        8'h72: rddata <= 12'd161;
        8'h73: rddata <= 12'd159;
        8'h74: rddata <= 12'd156;
        8'h75: rddata <= 12'd153;
        8'h76: rddata <= 12'd151;
        8'h77: rddata <= 12'd148;
        8'h78: rddata <= 12'd146;
        8'h79: rddata <= 12'd143;
        8'h7A: rddata <= 12'd141;
        8'h7B: rddata <= 12'd138;
        8'h7C: rddata <= 12'd136;
        8'h7D: rddata <= 12'd134;
        8'h7E: rddata <= 12'd131;
        8'h7F: rddata <= 12'd129;
        8'h80: rddata <= 12'd127;
        8'h81: rddata <= 12'd125;
        8'h82: rddata <= 12'd122;
        8'h83: rddata <= 12'd120;
        8'h84: rddata <= 12'd118;
        8'h85: rddata <= 12'd116;
        8'h86: rddata <= 12'd114;
        8'h87: rddata <= 12'd112;
        8'h88: rddata <= 12'd110;
        8'h89: rddata <= 12'd108;
        8'h8A: rddata <= 12'd106;
        8'h8B: rddata <= 12'd104;
        8'h8C: rddata <= 12'd102;
        8'h8D: rddata <= 12'd100;
        8'h8E: rddata <= 12'd98;
        8'h8F: rddata <= 12'd96;
        8'h90: rddata <= 12'd94;
        8'h91: rddata <= 12'd92;
        8'h92: rddata <= 12'd91;
        8'h93: rddata <= 12'd89;
        8'h94: rddata <= 12'd87;
        8'h95: rddata <= 12'd85;
        8'h96: rddata <= 12'd83;
        8'h97: rddata <= 12'd82;
        8'h98: rddata <= 12'd80;
        8'h99: rddata <= 12'd78;
        8'h9A: rddata <= 12'd77;
        8'h9B: rddata <= 12'd75;
        8'h9C: rddata <= 12'd74;
        8'h9D: rddata <= 12'd72;
        8'h9E: rddata <= 12'd70;
        8'h9F: rddata <= 12'd69;
        8'hA0: rddata <= 12'd67;
        8'hA1: rddata <= 12'd66;
        8'hA2: rddata <= 12'd64;
        8'hA3: rddata <= 12'd63;
        8'hA4: rddata <= 12'd62;
        8'hA5: rddata <= 12'd60;
        8'hA6: rddata <= 12'd59;
        8'hA7: rddata <= 12'd57;
        8'hA8: rddata <= 12'd56;
        8'hA9: rddata <= 12'd55;
        8'hAA: rddata <= 12'd53;
        8'hAB: rddata <= 12'd52;
        8'hAC: rddata <= 12'd51;
        8'hAD: rddata <= 12'd49;
        8'hAE: rddata <= 12'd48;
        8'hAF: rddata <= 12'd47;
        8'hB0: rddata <= 12'd46;
        8'hB1: rddata <= 12'd45;
        8'hB2: rddata <= 12'd43;
        8'hB3: rddata <= 12'd42;
        8'hB4: rddata <= 12'd41;
        8'hB5: rddata <= 12'd40;
        8'hB6: rddata <= 12'd39;
        8'hB7: rddata <= 12'd38;
        8'hB8: rddata <= 12'd37;
        8'hB9: rddata <= 12'd36;
        8'hBA: rddata <= 12'd35;
        8'hBB: rddata <= 12'd34;
        8'hBC: rddata <= 12'd33;
        8'hBD: rddata <= 12'd32;
        8'hBE: rddata <= 12'd31;
        8'hBF: rddata <= 12'd30;
        8'hC0: rddata <= 12'd29;
        8'hC1: rddata <= 12'd28;
        8'hC2: rddata <= 12'd27;
        8'hC3: rddata <= 12'd26;
        8'hC4: rddata <= 12'd25;
        8'hC5: rddata <= 12'd24;
        8'hC6: rddata <= 12'd23;
        8'hC7: rddata <= 12'd23;
        8'hC8: rddata <= 12'd22;
        8'hC9: rddata <= 12'd21;
        8'hCA: rddata <= 12'd20;
        8'hCB: rddata <= 12'd20;
        8'hCC: rddata <= 12'd19;
        8'hCD: rddata <= 12'd18;
        8'hCE: rddata <= 12'd17;
        8'hCF: rddata <= 12'd17;
        8'hD0: rddata <= 12'd16;
        8'hD1: rddata <= 12'd15;
        8'hD2: rddata <= 12'd15;
        8'hD3: rddata <= 12'd14;
        8'hD4: rddata <= 12'd13;
        8'hD5: rddata <= 12'd13;
        8'hD6: rddata <= 12'd12;
        8'hD7: rddata <= 12'd12;
        8'hD8: rddata <= 12'd11;
        8'hD9: rddata <= 12'd10;
        8'hDA: rddata <= 12'd10;
        8'hDB: rddata <= 12'd9;
        8'hDC: rddata <= 12'd9;
        8'hDD: rddata <= 12'd8;
        8'hDE: rddata <= 12'd8;
        8'hDF: rddata <= 12'd7;
        8'hE0: rddata <= 12'd7;
        8'hE1: rddata <= 12'd7;
        8'hE2: rddata <= 12'd6;
        8'hE3: rddata <= 12'd6;
        8'hE4: rddata <= 12'd5;
        8'hE5: rddata <= 12'd5;
        8'hE6: rddata <= 12'd5;
        8'hE7: rddata <= 12'd4;
        8'hE8: rddata <= 12'd4;
        8'hE9: rddata <= 12'd4;
        8'hEA: rddata <= 12'd3;
        8'hEB: rddata <= 12'd3;
        8'hEC: rddata <= 12'd3;
        8'hED: rddata <= 12'd2;
        8'hEE: rddata <= 12'd2;
        8'hEF: rddata <= 12'd2;
        8'hF0: rddata <= 12'd2;
        8'hF1: rddata <= 12'd1;
        8'hF2: rddata <= 12'd1;
        8'hF3: rddata <= 12'd1;
        8'hF4: rddata <= 12'd1;
        8'hF5: rddata <= 12'd1;
        8'hF6: rddata <= 12'd1;
        8'hF7: rddata <= 12'd1;
        8'hF8: rddata <= 12'd0;
        8'hF9: rddata <= 12'd0;
        8'hFA: rddata <= 12'd0;
        8'hFB: rddata <= 12'd0;
        8'hFC: rddata <= 12'd0;
        8'hFD: rddata <= 12'd0;
        8'hFE: rddata <= 12'd0;
        8'hFF: rddata <= 12'd0;
        default: rddata <= 12'd0;
    endcase

endmodule
