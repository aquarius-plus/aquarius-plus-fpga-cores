`default_nettype none
`timescale 1 ns / 1 ps

module bootrom(
    input  wire        clk,
    input  wire  [8:0] addr,
    output reg  [31:0] rddata
);

    always @(posedge clk) case (addr)
        9'h000:  rddata <= 32'h00001197;
        9'h001:  rddata <= 32'h00018193;
        9'h002:  rddata <= 32'h00080117;
        9'h003:  rddata <= 32'h7F810113;
        9'h004:  rddata <= 32'h00000293;
        9'h005:  rddata <= 32'h00000313;
        9'h006:  rddata <= 32'h00C0006F;
        9'h007:  rddata <= 32'h0002A023;
        9'h008:  rddata <= 32'h00428293;
        9'h009:  rddata <= 32'hFE62ECE3;
        9'h00A:  rddata <= 32'h00000293;
        9'h00B:  rddata <= 32'h00000313;
        9'h00C:  rddata <= 32'h00000397;
        9'h00D:  rddata <= 32'h2E038393;
        9'h00E:  rddata <= 32'h0140006F;
        9'h00F:  rddata <= 32'h0003AE03;
        9'h010:  rddata <= 32'h00438393;
        9'h011:  rddata <= 32'h01C2A023;
        9'h012:  rddata <= 32'h00428293;
        9'h013:  rddata <= 32'hFE62E8E3;
        9'h014:  rddata <= 32'h00000297;
        9'h015:  rddata <= 32'h00C28293;
        9'h016:  rddata <= 32'h00028067;
        9'h017:  rddata <= 32'hFF010113;
        9'h018:  rddata <= 32'h00112623;
        9'h019:  rddata <= 32'h00812423;
        9'h01A:  rddata <= 32'h00912223;
        9'h01B:  rddata <= 32'hFF0007B7;
        9'h01C:  rddata <= 32'h34100713;
        9'h01D:  rddata <= 32'h00E79023;
        9'h01E:  rddata <= 32'hFF5007B7;
        9'h01F:  rddata <= 32'h00100713;
        9'h020:  rddata <= 32'h00E7A423;
        9'h021:  rddata <= 32'h08300713;
        9'h022:  rddata <= 32'h00E7A023;
        9'h023:  rddata <= 32'h0007A703;
        9'h024:  rddata <= 32'h00277713;
        9'h025:  rddata <= 32'hFE071CE3;
        9'h026:  rddata <= 32'h00100713;
        9'h027:  rddata <= 32'h00E7A223;
        9'h028:  rddata <= 32'hFF0004B7;
        9'h029:  rddata <= 32'h34200793;
        9'h02A:  rddata <= 32'h00000537;
        9'h02B:  rddata <= 32'h00F49023;
        9'h02C:  rddata <= 32'h00000593;
        9'h02D:  rddata <= 32'hB0050513;
        9'h02E:  rddata <= 32'h12C000EF;
        9'h02F:  rddata <= 32'h34300793;
        9'h030:  rddata <= 32'h00F49023;
        9'h031:  rddata <= 32'h00050413;
        9'h032:  rddata <= 32'h00054E63;
        9'h033:  rddata <= 32'h00004637;
        9'h034:  rddata <= 32'h00000593;
        9'h035:  rddata <= 32'h174000EF;
        9'h036:  rddata <= 32'h00040513;
        9'h037:  rddata <= 32'h0CC000EF;
        9'h038:  rddata <= 32'h00000067;
        9'h039:  rddata <= 32'hFF0007B7;
        9'h03A:  rddata <= 32'h34400713;
        9'h03B:  rddata <= 32'h00E79023;
        9'h03C:  rddata <= 32'h0000006F;
        9'h03D:  rddata <= 32'hFF500737;
        9'h03E:  rddata <= 32'h00072783;
        9'h03F:  rddata <= 32'h0027F793;
        9'h040:  rddata <= 32'hFE079CE3;
        9'h041:  rddata <= 32'h00A72223;
        9'h042:  rddata <= 32'h00008067;
        9'h043:  rddata <= 32'hFF500737;
        9'h044:  rddata <= 32'h00072783;
        9'h045:  rddata <= 32'h0017F793;
        9'h046:  rddata <= 32'hFE078CE3;
        9'h047:  rddata <= 32'h00472503;
        9'h048:  rddata <= 32'h0FF57513;
        9'h049:  rddata <= 32'h00008067;
        9'h04A:  rddata <= 32'hFF5007B7;
        9'h04B:  rddata <= 32'h08300713;
        9'h04C:  rddata <= 32'h00E7A023;
        9'h04D:  rddata <= 32'hFC1FF06F;
        9'h04E:  rddata <= 32'hFF010113;
        9'h04F:  rddata <= 32'h00B505B3;
        9'h050:  rddata <= 32'h00912223;
        9'h051:  rddata <= 32'h01059493;
        9'h052:  rddata <= 32'h00812423;
        9'h053:  rddata <= 32'h00112623;
        9'h054:  rddata <= 32'h00050413;
        9'h055:  rddata <= 32'h0104D493;
        9'h056:  rddata <= 32'h01041793;
        9'h057:  rddata <= 32'h0107D793;
        9'h058:  rddata <= 32'h00F49C63;
        9'h059:  rddata <= 32'h00C12083;
        9'h05A:  rddata <= 32'h00812403;
        9'h05B:  rddata <= 32'h00412483;
        9'h05C:  rddata <= 32'h01010113;
        9'h05D:  rddata <= 32'h00008067;
        9'h05E:  rddata <= 32'h00044503;
        9'h05F:  rddata <= 32'h00140413;
        9'h060:  rddata <= 32'hF75FF0EF;
        9'h061:  rddata <= 32'hFD5FF06F;
        9'h062:  rddata <= 32'h00050793;
        9'h063:  rddata <= 32'h00000513;
        9'h064:  rddata <= 32'h00A78733;
        9'h065:  rddata <= 32'h00074703;
        9'h066:  rddata <= 32'h00071463;
        9'h067:  rddata <= 32'h00008067;
        9'h068:  rddata <= 32'h00150513;
        9'h069:  rddata <= 32'hFEDFF06F;
        9'h06A:  rddata <= 32'hFF010113;
        9'h06B:  rddata <= 32'h00812423;
        9'h06C:  rddata <= 32'h00050413;
        9'h06D:  rddata <= 32'h01100513;
        9'h06E:  rddata <= 32'h00112623;
        9'h06F:  rddata <= 32'hF6DFF0EF;
        9'h070:  rddata <= 32'h0FF47513;
        9'h071:  rddata <= 32'hF31FF0EF;
        9'h072:  rddata <= 32'hF45FF0EF;
        9'h073:  rddata <= 32'h00C12083;
        9'h074:  rddata <= 32'h00812403;
        9'h075:  rddata <= 32'h01851513;
        9'h076:  rddata <= 32'h41855513;
        9'h077:  rddata <= 32'h01010113;
        9'h078:  rddata <= 32'h00008067;
        9'h079:  rddata <= 32'hFF010113;
        9'h07A:  rddata <= 32'h00812423;
        9'h07B:  rddata <= 32'h00050413;
        9'h07C:  rddata <= 32'h01000513;
        9'h07D:  rddata <= 32'h00112623;
        9'h07E:  rddata <= 32'h00912223;
        9'h07F:  rddata <= 32'h00058493;
        9'h080:  rddata <= 32'hF29FF0EF;
        9'h081:  rddata <= 32'h00048513;
        9'h082:  rddata <= 32'hEEDFF0EF;
        9'h083:  rddata <= 32'h00040513;
        9'h084:  rddata <= 32'hF79FF0EF;
        9'h085:  rddata <= 32'h00150593;
        9'h086:  rddata <= 32'h01059593;
        9'h087:  rddata <= 32'h00040513;
        9'h088:  rddata <= 32'h0105D593;
        9'h089:  rddata <= 32'hF15FF0EF;
        9'h08A:  rddata <= 32'hEE5FF0EF;
        9'h08B:  rddata <= 32'h00C12083;
        9'h08C:  rddata <= 32'h00812403;
        9'h08D:  rddata <= 32'h01851513;
        9'h08E:  rddata <= 32'h00412483;
        9'h08F:  rddata <= 32'h41855513;
        9'h090:  rddata <= 32'h01010113;
        9'h091:  rddata <= 32'h00008067;
        9'h092:  rddata <= 32'hFF010113;
        9'h093:  rddata <= 32'h00912223;
        9'h094:  rddata <= 32'h00050493;
        9'h095:  rddata <= 32'h01200513;
        9'h096:  rddata <= 32'h00112623;
        9'h097:  rddata <= 32'h00812423;
        9'h098:  rddata <= 32'h01212023;
        9'h099:  rddata <= 32'h00060413;
        9'h09A:  rddata <= 32'h00058913;
        9'h09B:  rddata <= 32'hEBDFF0EF;
        9'h09C:  rddata <= 32'h0FF4F513;
        9'h09D:  rddata <= 32'hE81FF0EF;
        9'h09E:  rddata <= 32'h0FF47513;
        9'h09F:  rddata <= 32'hE79FF0EF;
        9'h0A0:  rddata <= 32'h00845513;
        9'h0A1:  rddata <= 32'hE71FF0EF;
        9'h0A2:  rddata <= 32'hE85FF0EF;
        9'h0A3:  rddata <= 32'h01851513;
        9'h0A4:  rddata <= 32'h41855513;
        9'h0A5:  rddata <= 32'h04054063;
        9'h0A6:  rddata <= 32'hE75FF0EF;
        9'h0A7:  rddata <= 32'h01051413;
        9'h0A8:  rddata <= 32'hE6DFF0EF;
        9'h0A9:  rddata <= 32'h41045413;
        9'h0AA:  rddata <= 32'h00851513;
        9'h0AB:  rddata <= 32'h00A467B3;
        9'h0AC:  rddata <= 32'h01079493;
        9'h0AD:  rddata <= 32'h00F907B3;
        9'h0AE:  rddata <= 32'h01079413;
        9'h0AF:  rddata <= 32'h4104D493;
        9'h0B0:  rddata <= 32'h01045413;
        9'h0B1:  rddata <= 32'h01091793;
        9'h0B2:  rddata <= 32'h0107D793;
        9'h0B3:  rddata <= 32'h02F41063;
        9'h0B4:  rddata <= 32'h00048513;
        9'h0B5:  rddata <= 32'h00C12083;
        9'h0B6:  rddata <= 32'h00812403;
        9'h0B7:  rddata <= 32'h00412483;
        9'h0B8:  rddata <= 32'h00012903;
        9'h0B9:  rddata <= 32'h01010113;
        9'h0BA:  rddata <= 32'h00008067;
        9'h0BB:  rddata <= 32'h00190913;
        9'h0BC:  rddata <= 32'hE1DFF0EF;
        9'h0BD:  rddata <= 32'hFEA90FA3;
        9'h0BE:  rddata <= 32'hFCDFF06F;
        9'h0BF:  rddata <= 32'h00000000;
        9'h0C0:  rddata <= 32'h32337161;
        9'h0C1:  rddata <= 32'h6D6F722E;
        9'h0C2:  rddata <= 32'h00000000;
        default: rddata <= 32'h00000000;
    endcase

endmodule
