`default_nettype none
`timescale 1 ns / 1 ps

(* rom_style = "distributed" *)
module lut_pan_r(
    input  wire  [6:0] idx,
    output reg   [7:0] value
);

    always @* case (idx)
        7'h00: value = 8'h00;
        7'h01: value = 8'h00;
        7'h02: value = 8'h03;
        7'h03: value = 8'h06;
        7'h04: value = 8'h09;
        7'h05: value = 8'h0c;
        7'h06: value = 8'h0f;
        7'h07: value = 8'h13;
        7'h08: value = 8'h16;
        7'h09: value = 8'h19;
        7'h0A: value = 8'h1c;
        7'h0B: value = 8'h1f;
        7'h0C: value = 8'h22;
        7'h0D: value = 8'h26;
        7'h0E: value = 8'h29;
        7'h0F: value = 8'h2c;
        7'h10: value = 8'h2f;
        7'h11: value = 8'h32;
        7'h12: value = 8'h35;
        7'h13: value = 8'h38;
        7'h14: value = 8'h3b;
        7'h15: value = 8'h3e;
        7'h16: value = 8'h41;
        7'h17: value = 8'h45;
        7'h18: value = 8'h48;
        7'h19: value = 8'h4b;
        7'h1A: value = 8'h4e;
        7'h1B: value = 8'h51;
        7'h1C: value = 8'h54;
        7'h1D: value = 8'h57;
        7'h1E: value = 8'h5a;
        7'h1F: value = 8'h5d;
        7'h20: value = 8'h60;
        7'h21: value = 8'h63;
        7'h22: value = 8'h65;
        7'h23: value = 8'h68;
        7'h24: value = 8'h6b;
        7'h25: value = 8'h6e;
        7'h26: value = 8'h71;
        7'h27: value = 8'h74;
        7'h28: value = 8'h77;
        7'h29: value = 8'h79;
        7'h2A: value = 8'h7c;
        7'h2B: value = 8'h7f;
        7'h2C: value = 8'h82;
        7'h2D: value = 8'h84;
        7'h2E: value = 8'h87;
        7'h2F: value = 8'h8a;
        7'h30: value = 8'h8d;
        7'h31: value = 8'h8f;
        7'h32: value = 8'h92;
        7'h33: value = 8'h94;
        7'h34: value = 8'h97;
        7'h35: value = 8'h99;
        7'h36: value = 8'h9c;
        7'h37: value = 8'h9e;
        7'h38: value = 8'ha1;
        7'h39: value = 8'ha3;
        7'h3A: value = 8'ha6;
        7'h3B: value = 8'ha8;
        7'h3C: value = 8'hab;
        7'h3D: value = 8'had;
        7'h3E: value = 8'haf;
        7'h3F: value = 8'hb2;
        7'h40: value = 8'hb4;
        7'h41: value = 8'hb6;
        7'h42: value = 8'hb8;
        7'h43: value = 8'hba;
        7'h44: value = 8'hbd;
        7'h45: value = 8'hbf;
        7'h46: value = 8'hc1;
        7'h47: value = 8'hc3;
        7'h48: value = 8'hc5;
        7'h49: value = 8'hc7;
        7'h4A: value = 8'hc9;
        7'h4B: value = 8'hcb;
        7'h4C: value = 8'hcd;
        7'h4D: value = 8'hcf;
        7'h4E: value = 8'hd0;
        7'h4F: value = 8'hd2;
        7'h50: value = 8'hd4;
        7'h51: value = 8'hd6;
        7'h52: value = 8'hd7;
        7'h53: value = 8'hd9;
        7'h54: value = 8'hdb;
        7'h55: value = 8'hdc;
        7'h56: value = 8'hde;
        7'h57: value = 8'hdf;
        7'h58: value = 8'he1;
        7'h59: value = 8'he2;
        7'h5A: value = 8'he4;
        7'h5B: value = 8'he5;
        7'h5C: value = 8'he7;
        7'h5D: value = 8'he8;
        7'h5E: value = 8'he9;
        7'h5F: value = 8'hea;
        7'h60: value = 8'hec;
        7'h61: value = 8'hed;
        7'h62: value = 8'hee;
        7'h63: value = 8'hef;
        7'h64: value = 8'hf0;
        7'h65: value = 8'hf1;
        7'h66: value = 8'hf2;
        7'h67: value = 8'hf3;
        7'h68: value = 8'hf4;
        7'h69: value = 8'hf5;
        7'h6A: value = 8'hf6;
        7'h6B: value = 8'hf7;
        7'h6C: value = 8'hf7;
        7'h6D: value = 8'hf8;
        7'h6E: value = 8'hf9;
        7'h6F: value = 8'hf9;
        7'h70: value = 8'hfa;
        7'h71: value = 8'hfb;
        7'h72: value = 8'hfb;
        7'h73: value = 8'hfc;
        7'h74: value = 8'hfc;
        7'h75: value = 8'hfd;
        7'h76: value = 8'hfd;
        7'h77: value = 8'hfd;
        7'h78: value = 8'hfe;
        7'h79: value = 8'hfe;
        7'h7A: value = 8'hfe;
        7'h7B: value = 8'hfe;
        7'h7C: value = 8'hfe;
        7'h7D: value = 8'hfe;
        7'h7E: value = 8'hfe;
        7'h7F: value = 8'hff;
        default: value = 8'h0;
    endcase

endmodule
