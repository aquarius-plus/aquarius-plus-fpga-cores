`default_nettype none
`timescale 1 ns / 1 ps

(* rom_style = "distributed" *)
module lut_logsin(
    input  wire        clk,
    input  wire  [7:0] idx,
    output reg  [11:0] value
);

    always @(posedge clk) case (idx)
        8'h00: value <= 12'd2137;
        8'h01: value <= 12'd1731;
        8'h02: value <= 12'd1543;
        8'h03: value <= 12'd1419;
        8'h04: value <= 12'd1326;
        8'h05: value <= 12'd1252;
        8'h06: value <= 12'd1190;
        8'h07: value <= 12'd1137;
        8'h08: value <= 12'd1091;
        8'h09: value <= 12'd1050;
        8'h0A: value <= 12'd1013;
        8'h0B: value <= 12'd979;
        8'h0C: value <= 12'd949;
        8'h0D: value <= 12'd920;
        8'h0E: value <= 12'd894;
        8'h0F: value <= 12'd869;
        8'h10: value <= 12'd846;
        8'h11: value <= 12'd825;
        8'h12: value <= 12'd804;
        8'h13: value <= 12'd785;
        8'h14: value <= 12'd767;
        8'h15: value <= 12'd749;
        8'h16: value <= 12'd732;
        8'h17: value <= 12'd717;
        8'h18: value <= 12'd701;
        8'h19: value <= 12'd687;
        8'h1A: value <= 12'd672;
        8'h1B: value <= 12'd659;
        8'h1C: value <= 12'd646;
        8'h1D: value <= 12'd633;
        8'h1E: value <= 12'd621;
        8'h1F: value <= 12'd609;
        8'h20: value <= 12'd598;
        8'h21: value <= 12'd587;
        8'h22: value <= 12'd576;
        8'h23: value <= 12'd566;
        8'h24: value <= 12'd556;
        8'h25: value <= 12'd546;
        8'h26: value <= 12'd536;
        8'h27: value <= 12'd527;
        8'h28: value <= 12'd518;
        8'h29: value <= 12'd509;
        8'h2A: value <= 12'd501;
        8'h2B: value <= 12'd492;
        8'h2C: value <= 12'd484;
        8'h2D: value <= 12'd476;
        8'h2E: value <= 12'd468;
        8'h2F: value <= 12'd461;
        8'h30: value <= 12'd453;
        8'h31: value <= 12'd446;
        8'h32: value <= 12'd439;
        8'h33: value <= 12'd432;
        8'h34: value <= 12'd425;
        8'h35: value <= 12'd418;
        8'h36: value <= 12'd411;
        8'h37: value <= 12'd405;
        8'h38: value <= 12'd399;
        8'h39: value <= 12'd392;
        8'h3A: value <= 12'd386;
        8'h3B: value <= 12'd380;
        8'h3C: value <= 12'd375;
        8'h3D: value <= 12'd369;
        8'h3E: value <= 12'd363;
        8'h3F: value <= 12'd358;
        8'h40: value <= 12'd352;
        8'h41: value <= 12'd347;
        8'h42: value <= 12'd341;
        8'h43: value <= 12'd336;
        8'h44: value <= 12'd331;
        8'h45: value <= 12'd326;
        8'h46: value <= 12'd321;
        8'h47: value <= 12'd316;
        8'h48: value <= 12'd311;
        8'h49: value <= 12'd307;
        8'h4A: value <= 12'd302;
        8'h4B: value <= 12'd297;
        8'h4C: value <= 12'd293;
        8'h4D: value <= 12'd289;
        8'h4E: value <= 12'd284;
        8'h4F: value <= 12'd280;
        8'h50: value <= 12'd276;
        8'h51: value <= 12'd271;
        8'h52: value <= 12'd267;
        8'h53: value <= 12'd263;
        8'h54: value <= 12'd259;
        8'h55: value <= 12'd255;
        8'h56: value <= 12'd251;
        8'h57: value <= 12'd248;
        8'h58: value <= 12'd244;
        8'h59: value <= 12'd240;
        8'h5A: value <= 12'd236;
        8'h5B: value <= 12'd233;
        8'h5C: value <= 12'd229;
        8'h5D: value <= 12'd226;
        8'h5E: value <= 12'd222;
        8'h5F: value <= 12'd219;
        8'h60: value <= 12'd215;
        8'h61: value <= 12'd212;
        8'h62: value <= 12'd209;
        8'h63: value <= 12'd205;
        8'h64: value <= 12'd202;
        8'h65: value <= 12'd199;
        8'h66: value <= 12'd196;
        8'h67: value <= 12'd193;
        8'h68: value <= 12'd190;
        8'h69: value <= 12'd187;
        8'h6A: value <= 12'd184;
        8'h6B: value <= 12'd181;
        8'h6C: value <= 12'd178;
        8'h6D: value <= 12'd175;
        8'h6E: value <= 12'd172;
        8'h6F: value <= 12'd169;
        8'h70: value <= 12'd167;
        8'h71: value <= 12'd164;
        8'h72: value <= 12'd161;
        8'h73: value <= 12'd159;
        8'h74: value <= 12'd156;
        8'h75: value <= 12'd153;
        8'h76: value <= 12'd151;
        8'h77: value <= 12'd148;
        8'h78: value <= 12'd146;
        8'h79: value <= 12'd143;
        8'h7A: value <= 12'd141;
        8'h7B: value <= 12'd138;
        8'h7C: value <= 12'd136;
        8'h7D: value <= 12'd134;
        8'h7E: value <= 12'd131;
        8'h7F: value <= 12'd129;
        8'h80: value <= 12'd127;
        8'h81: value <= 12'd125;
        8'h82: value <= 12'd122;
        8'h83: value <= 12'd120;
        8'h84: value <= 12'd118;
        8'h85: value <= 12'd116;
        8'h86: value <= 12'd114;
        8'h87: value <= 12'd112;
        8'h88: value <= 12'd110;
        8'h89: value <= 12'd108;
        8'h8A: value <= 12'd106;
        8'h8B: value <= 12'd104;
        8'h8C: value <= 12'd102;
        8'h8D: value <= 12'd100;
        8'h8E: value <= 12'd98;
        8'h8F: value <= 12'd96;
        8'h90: value <= 12'd94;
        8'h91: value <= 12'd92;
        8'h92: value <= 12'd91;
        8'h93: value <= 12'd89;
        8'h94: value <= 12'd87;
        8'h95: value <= 12'd85;
        8'h96: value <= 12'd83;
        8'h97: value <= 12'd82;
        8'h98: value <= 12'd80;
        8'h99: value <= 12'd78;
        8'h9A: value <= 12'd77;
        8'h9B: value <= 12'd75;
        8'h9C: value <= 12'd74;
        8'h9D: value <= 12'd72;
        8'h9E: value <= 12'd70;
        8'h9F: value <= 12'd69;
        8'hA0: value <= 12'd67;
        8'hA1: value <= 12'd66;
        8'hA2: value <= 12'd64;
        8'hA3: value <= 12'd63;
        8'hA4: value <= 12'd62;
        8'hA5: value <= 12'd60;
        8'hA6: value <= 12'd59;
        8'hA7: value <= 12'd57;
        8'hA8: value <= 12'd56;
        8'hA9: value <= 12'd55;
        8'hAA: value <= 12'd53;
        8'hAB: value <= 12'd52;
        8'hAC: value <= 12'd51;
        8'hAD: value <= 12'd49;
        8'hAE: value <= 12'd48;
        8'hAF: value <= 12'd47;
        8'hB0: value <= 12'd46;
        8'hB1: value <= 12'd45;
        8'hB2: value <= 12'd43;
        8'hB3: value <= 12'd42;
        8'hB4: value <= 12'd41;
        8'hB5: value <= 12'd40;
        8'hB6: value <= 12'd39;
        8'hB7: value <= 12'd38;
        8'hB8: value <= 12'd37;
        8'hB9: value <= 12'd36;
        8'hBA: value <= 12'd35;
        8'hBB: value <= 12'd34;
        8'hBC: value <= 12'd33;
        8'hBD: value <= 12'd32;
        8'hBE: value <= 12'd31;
        8'hBF: value <= 12'd30;
        8'hC0: value <= 12'd29;
        8'hC1: value <= 12'd28;
        8'hC2: value <= 12'd27;
        8'hC3: value <= 12'd26;
        8'hC4: value <= 12'd25;
        8'hC5: value <= 12'd24;
        8'hC6: value <= 12'd23;
        8'hC7: value <= 12'd23;
        8'hC8: value <= 12'd22;
        8'hC9: value <= 12'd21;
        8'hCA: value <= 12'd20;
        8'hCB: value <= 12'd20;
        8'hCC: value <= 12'd19;
        8'hCD: value <= 12'd18;
        8'hCE: value <= 12'd17;
        8'hCF: value <= 12'd17;
        8'hD0: value <= 12'd16;
        8'hD1: value <= 12'd15;
        8'hD2: value <= 12'd15;
        8'hD3: value <= 12'd14;
        8'hD4: value <= 12'd13;
        8'hD5: value <= 12'd13;
        8'hD6: value <= 12'd12;
        8'hD7: value <= 12'd12;
        8'hD8: value <= 12'd11;
        8'hD9: value <= 12'd10;
        8'hDA: value <= 12'd10;
        8'hDB: value <= 12'd9;
        8'hDC: value <= 12'd9;
        8'hDD: value <= 12'd8;
        8'hDE: value <= 12'd8;
        8'hDF: value <= 12'd7;
        8'hE0: value <= 12'd7;
        8'hE1: value <= 12'd7;
        8'hE2: value <= 12'd6;
        8'hE3: value <= 12'd6;
        8'hE4: value <= 12'd5;
        8'hE5: value <= 12'd5;
        8'hE6: value <= 12'd5;
        8'hE7: value <= 12'd4;
        8'hE8: value <= 12'd4;
        8'hE9: value <= 12'd4;
        8'hEA: value <= 12'd3;
        8'hEB: value <= 12'd3;
        8'hEC: value <= 12'd3;
        8'hED: value <= 12'd2;
        8'hEE: value <= 12'd2;
        8'hEF: value <= 12'd2;
        8'hF0: value <= 12'd2;
        8'hF1: value <= 12'd1;
        8'hF2: value <= 12'd1;
        8'hF3: value <= 12'd1;
        8'hF4: value <= 12'd1;
        8'hF5: value <= 12'd1;
        8'hF6: value <= 12'd1;
        8'hF7: value <= 12'd1;
        8'hF8: value <= 12'd0;
        8'hF9: value <= 12'd0;
        8'hFA: value <= 12'd0;
        8'hFB: value <= 12'd0;
        8'hFC: value <= 12'd0;
        8'hFD: value <= 12'd0;
        8'hFE: value <= 12'd0;
        8'hFF: value <= 12'd0;
        default: value <= 12'd0;
    endcase

endmodule
