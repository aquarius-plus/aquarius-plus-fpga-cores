`default_nettype none
`timescale 1 ns / 1 ps

(* rom_style = "distributed" *)
module fm_exp_rom(
    input  wire  [7:0] idx,
    output reg   [9:0] value
);

    always @* case (idx)
        8'h00: value = 10'h3fa;
        8'h01: value = 10'h3f5;
        8'h02: value = 10'h3ef;
        8'h03: value = 10'h3ea;
        8'h04: value = 10'h3e4;
        8'h05: value = 10'h3df;
        8'h06: value = 10'h3da;
        8'h07: value = 10'h3d4;
        8'h08: value = 10'h3cf;
        8'h09: value = 10'h3c9;
        8'h0A: value = 10'h3c4;
        8'h0B: value = 10'h3bf;
        8'h0C: value = 10'h3b9;
        8'h0D: value = 10'h3b4;
        8'h0E: value = 10'h3ae;
        8'h0F: value = 10'h3a9;
        8'h10: value = 10'h3a4;
        8'h11: value = 10'h39f;
        8'h12: value = 10'h399;
        8'h13: value = 10'h394;
        8'h14: value = 10'h38f;
        8'h15: value = 10'h38a;
        8'h16: value = 10'h384;
        8'h17: value = 10'h37f;
        8'h18: value = 10'h37a;
        8'h19: value = 10'h375;
        8'h1A: value = 10'h370;
        8'h1B: value = 10'h36a;
        8'h1C: value = 10'h365;
        8'h1D: value = 10'h360;
        8'h1E: value = 10'h35b;
        8'h1F: value = 10'h356;
        8'h20: value = 10'h351;
        8'h21: value = 10'h34c;
        8'h22: value = 10'h347;
        8'h23: value = 10'h342;
        8'h24: value = 10'h33d;
        8'h25: value = 10'h338;
        8'h26: value = 10'h333;
        8'h27: value = 10'h32e;
        8'h28: value = 10'h329;
        8'h29: value = 10'h324;
        8'h2A: value = 10'h31f;
        8'h2B: value = 10'h31a;
        8'h2C: value = 10'h315;
        8'h2D: value = 10'h310;
        8'h2E: value = 10'h30b;
        8'h2F: value = 10'h306;
        8'h30: value = 10'h302;
        8'h31: value = 10'h2fd;
        8'h32: value = 10'h2f8;
        8'h33: value = 10'h2f3;
        8'h34: value = 10'h2ee;
        8'h35: value = 10'h2e9;
        8'h36: value = 10'h2e5;
        8'h37: value = 10'h2e0;
        8'h38: value = 10'h2db;
        8'h39: value = 10'h2d6;
        8'h3A: value = 10'h2d2;
        8'h3B: value = 10'h2cd;
        8'h3C: value = 10'h2c8;
        8'h3D: value = 10'h2c4;
        8'h3E: value = 10'h2bf;
        8'h3F: value = 10'h2ba;
        8'h40: value = 10'h2b5;
        8'h41: value = 10'h2b1;
        8'h42: value = 10'h2ac;
        8'h43: value = 10'h2a8;
        8'h44: value = 10'h2a3;
        8'h45: value = 10'h29e;
        8'h46: value = 10'h29a;
        8'h47: value = 10'h295;
        8'h48: value = 10'h291;
        8'h49: value = 10'h28c;
        8'h4A: value = 10'h288;
        8'h4B: value = 10'h283;
        8'h4C: value = 10'h27f;
        8'h4D: value = 10'h27a;
        8'h4E: value = 10'h276;
        8'h4F: value = 10'h271;
        8'h50: value = 10'h26d;
        8'h51: value = 10'h268;
        8'h52: value = 10'h264;
        8'h53: value = 10'h25f;
        8'h54: value = 10'h25b;
        8'h55: value = 10'h257;
        8'h56: value = 10'h252;
        8'h57: value = 10'h24e;
        8'h58: value = 10'h249;
        8'h59: value = 10'h245;
        8'h5A: value = 10'h241;
        8'h5B: value = 10'h23c;
        8'h5C: value = 10'h238;
        8'h5D: value = 10'h234;
        8'h5E: value = 10'h230;
        8'h5F: value = 10'h22b;
        8'h60: value = 10'h227;
        8'h61: value = 10'h223;
        8'h62: value = 10'h21e;
        8'h63: value = 10'h21a;
        8'h64: value = 10'h216;
        8'h65: value = 10'h212;
        8'h66: value = 10'h20e;
        8'h67: value = 10'h209;
        8'h68: value = 10'h205;
        8'h69: value = 10'h201;
        8'h6A: value = 10'h1fd;
        8'h6B: value = 10'h1f9;
        8'h6C: value = 10'h1f5;
        8'h6D: value = 10'h1f0;
        8'h6E: value = 10'h1ec;
        8'h6F: value = 10'h1e8;
        8'h70: value = 10'h1e4;
        8'h71: value = 10'h1e0;
        8'h72: value = 10'h1dc;
        8'h73: value = 10'h1d8;
        8'h74: value = 10'h1d4;
        8'h75: value = 10'h1d0;
        8'h76: value = 10'h1cc;
        8'h77: value = 10'h1c8;
        8'h78: value = 10'h1c4;
        8'h79: value = 10'h1c0;
        8'h7A: value = 10'h1bc;
        8'h7B: value = 10'h1b8;
        8'h7C: value = 10'h1b4;
        8'h7D: value = 10'h1b0;
        8'h7E: value = 10'h1ac;
        8'h7F: value = 10'h1a8;
        8'h80: value = 10'h1a4;
        8'h81: value = 10'h1a0;
        8'h82: value = 10'h19c;
        8'h83: value = 10'h199;
        8'h84: value = 10'h195;
        8'h85: value = 10'h191;
        8'h86: value = 10'h18d;
        8'h87: value = 10'h189;
        8'h88: value = 10'h185;
        8'h89: value = 10'h181;
        8'h8A: value = 10'h17e;
        8'h8B: value = 10'h17a;
        8'h8C: value = 10'h176;
        8'h8D: value = 10'h172;
        8'h8E: value = 10'h16f;
        8'h8F: value = 10'h16b;
        8'h90: value = 10'h167;
        8'h91: value = 10'h163;
        8'h92: value = 10'h160;
        8'h93: value = 10'h15c;
        8'h94: value = 10'h158;
        8'h95: value = 10'h154;
        8'h96: value = 10'h151;
        8'h97: value = 10'h14d;
        8'h98: value = 10'h149;
        8'h99: value = 10'h146;
        8'h9A: value = 10'h142;
        8'h9B: value = 10'h13e;
        8'h9C: value = 10'h13b;
        8'h9D: value = 10'h137;
        8'h9E: value = 10'h134;
        8'h9F: value = 10'h130;
        8'hA0: value = 10'h12c;
        8'hA1: value = 10'h129;
        8'hA2: value = 10'h125;
        8'hA3: value = 10'h122;
        8'hA4: value = 10'h11e;
        8'hA5: value = 10'h11b;
        8'hA6: value = 10'h117;
        8'hA7: value = 10'h114;
        8'hA8: value = 10'h110;
        8'hA9: value = 10'h10c;
        8'hAA: value = 10'h109;
        8'hAB: value = 10'h106;
        8'hAC: value = 10'h102;
        8'hAD: value = 10'h0ff;
        8'hAE: value = 10'h0fb;
        8'hAF: value = 10'h0f8;
        8'hB0: value = 10'h0f4;
        8'hB1: value = 10'h0f1;
        8'hB2: value = 10'h0ed;
        8'hB3: value = 10'h0ea;
        8'hB4: value = 10'h0e7;
        8'hB5: value = 10'h0e3;
        8'hB6: value = 10'h0e0;
        8'hB7: value = 10'h0dc;
        8'hB8: value = 10'h0d9;
        8'hB9: value = 10'h0d6;
        8'hBA: value = 10'h0d2;
        8'hBB: value = 10'h0cf;
        8'hBC: value = 10'h0cc;
        8'hBD: value = 10'h0c8;
        8'hBE: value = 10'h0c5;
        8'hBF: value = 10'h0c2;
        8'hC0: value = 10'h0be;
        8'hC1: value = 10'h0bb;
        8'hC2: value = 10'h0b8;
        8'hC3: value = 10'h0b5;
        8'hC4: value = 10'h0b1;
        8'hC5: value = 10'h0ae;
        8'hC6: value = 10'h0ab;
        8'hC7: value = 10'h0a8;
        8'hC8: value = 10'h0a4;
        8'hC9: value = 10'h0a1;
        8'hCA: value = 10'h09e;
        8'hCB: value = 10'h09b;
        8'hCC: value = 10'h098;
        8'hCD: value = 10'h094;
        8'hCE: value = 10'h091;
        8'hCF: value = 10'h08e;
        8'hD0: value = 10'h08b;
        8'hD1: value = 10'h088;
        8'hD2: value = 10'h085;
        8'hD3: value = 10'h082;
        8'hD4: value = 10'h07e;
        8'hD5: value = 10'h07b;
        8'hD6: value = 10'h078;
        8'hD7: value = 10'h075;
        8'hD8: value = 10'h072;
        8'hD9: value = 10'h06f;
        8'hDA: value = 10'h06c;
        8'hDB: value = 10'h069;
        8'hDC: value = 10'h066;
        8'hDD: value = 10'h063;
        8'hDE: value = 10'h060;
        8'hDF: value = 10'h05d;
        8'hE0: value = 10'h05a;
        8'hE1: value = 10'h057;
        8'hE2: value = 10'h054;
        8'hE3: value = 10'h051;
        8'hE4: value = 10'h04e;
        8'hE5: value = 10'h04b;
        8'hE6: value = 10'h048;
        8'hE7: value = 10'h045;
        8'hE8: value = 10'h042;
        8'hE9: value = 10'h03f;
        8'hEA: value = 10'h03c;
        8'hEB: value = 10'h039;
        8'hEC: value = 10'h036;
        8'hED: value = 10'h033;
        8'hEE: value = 10'h030;
        8'hEF: value = 10'h02d;
        8'hF0: value = 10'h02a;
        8'hF1: value = 10'h028;
        8'hF2: value = 10'h025;
        8'hF3: value = 10'h022;
        8'hF4: value = 10'h01f;
        8'hF5: value = 10'h01c;
        8'hF6: value = 10'h019;
        8'hF7: value = 10'h016;
        8'hF8: value = 10'h014;
        8'hF9: value = 10'h011;
        8'hFA: value = 10'h00e;
        8'hFB: value = 10'h00b;
        8'hFC: value = 10'h008;
        8'hFD: value = 10'h006;
        8'hFE: value = 10'h003;
        8'hFF: value = 10'h000;
        default: value = 10'h0;
    endcase

endmodule
