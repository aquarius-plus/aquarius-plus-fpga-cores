`default_nettype none
`timescale 1 ns / 1 ps

module fmlut(
    input  wire        clk,
    input  wire  [8:0] addr,
    output reg  [11:0] rddata
);

    always @(posedge clk) case (addr)
        9'h000:  rddata <= 12'd2137;
        9'h001:  rddata <= 12'd1731;
        9'h002:  rddata <= 12'd1543;
        9'h003:  rddata <= 12'd1419;
        9'h004:  rddata <= 12'd1326;
        9'h005:  rddata <= 12'd1252;
        9'h006:  rddata <= 12'd1190;
        9'h007:  rddata <= 12'd1137;
        9'h008:  rddata <= 12'd1091;
        9'h009:  rddata <= 12'd1050;
        9'h00A:  rddata <= 12'd1013;
        9'h00B:  rddata <= 12'd979;
        9'h00C:  rddata <= 12'd949;
        9'h00D:  rddata <= 12'd920;
        9'h00E:  rddata <= 12'd894;
        9'h00F:  rddata <= 12'd869;
        9'h010:  rddata <= 12'd846;
        9'h011:  rddata <= 12'd825;
        9'h012:  rddata <= 12'd804;
        9'h013:  rddata <= 12'd785;
        9'h014:  rddata <= 12'd767;
        9'h015:  rddata <= 12'd749;
        9'h016:  rddata <= 12'd732;
        9'h017:  rddata <= 12'd717;
        9'h018:  rddata <= 12'd701;
        9'h019:  rddata <= 12'd687;
        9'h01A:  rddata <= 12'd672;
        9'h01B:  rddata <= 12'd659;
        9'h01C:  rddata <= 12'd646;
        9'h01D:  rddata <= 12'd633;
        9'h01E:  rddata <= 12'd621;
        9'h01F:  rddata <= 12'd609;
        9'h020:  rddata <= 12'd598;
        9'h021:  rddata <= 12'd587;
        9'h022:  rddata <= 12'd576;
        9'h023:  rddata <= 12'd566;
        9'h024:  rddata <= 12'd556;
        9'h025:  rddata <= 12'd546;
        9'h026:  rddata <= 12'd536;
        9'h027:  rddata <= 12'd527;
        9'h028:  rddata <= 12'd518;
        9'h029:  rddata <= 12'd509;
        9'h02A:  rddata <= 12'd501;
        9'h02B:  rddata <= 12'd492;
        9'h02C:  rddata <= 12'd484;
        9'h02D:  rddata <= 12'd476;
        9'h02E:  rddata <= 12'd468;
        9'h02F:  rddata <= 12'd461;
        9'h030:  rddata <= 12'd453;
        9'h031:  rddata <= 12'd446;
        9'h032:  rddata <= 12'd439;
        9'h033:  rddata <= 12'd432;
        9'h034:  rddata <= 12'd425;
        9'h035:  rddata <= 12'd418;
        9'h036:  rddata <= 12'd411;
        9'h037:  rddata <= 12'd405;
        9'h038:  rddata <= 12'd399;
        9'h039:  rddata <= 12'd392;
        9'h03A:  rddata <= 12'd386;
        9'h03B:  rddata <= 12'd380;
        9'h03C:  rddata <= 12'd375;
        9'h03D:  rddata <= 12'd369;
        9'h03E:  rddata <= 12'd363;
        9'h03F:  rddata <= 12'd358;
        9'h040:  rddata <= 12'd352;
        9'h041:  rddata <= 12'd347;
        9'h042:  rddata <= 12'd341;
        9'h043:  rddata <= 12'd336;
        9'h044:  rddata <= 12'd331;
        9'h045:  rddata <= 12'd326;
        9'h046:  rddata <= 12'd321;
        9'h047:  rddata <= 12'd316;
        9'h048:  rddata <= 12'd311;
        9'h049:  rddata <= 12'd307;
        9'h04A:  rddata <= 12'd302;
        9'h04B:  rddata <= 12'd297;
        9'h04C:  rddata <= 12'd293;
        9'h04D:  rddata <= 12'd289;
        9'h04E:  rddata <= 12'd284;
        9'h04F:  rddata <= 12'd280;
        9'h050:  rddata <= 12'd276;
        9'h051:  rddata <= 12'd271;
        9'h052:  rddata <= 12'd267;
        9'h053:  rddata <= 12'd263;
        9'h054:  rddata <= 12'd259;
        9'h055:  rddata <= 12'd255;
        9'h056:  rddata <= 12'd251;
        9'h057:  rddata <= 12'd248;
        9'h058:  rddata <= 12'd244;
        9'h059:  rddata <= 12'd240;
        9'h05A:  rddata <= 12'd236;
        9'h05B:  rddata <= 12'd233;
        9'h05C:  rddata <= 12'd229;
        9'h05D:  rddata <= 12'd226;
        9'h05E:  rddata <= 12'd222;
        9'h05F:  rddata <= 12'd219;
        9'h060:  rddata <= 12'd215;
        9'h061:  rddata <= 12'd212;
        9'h062:  rddata <= 12'd209;
        9'h063:  rddata <= 12'd205;
        9'h064:  rddata <= 12'd202;
        9'h065:  rddata <= 12'd199;
        9'h066:  rddata <= 12'd196;
        9'h067:  rddata <= 12'd193;
        9'h068:  rddata <= 12'd190;
        9'h069:  rddata <= 12'd187;
        9'h06A:  rddata <= 12'd184;
        9'h06B:  rddata <= 12'd181;
        9'h06C:  rddata <= 12'd178;
        9'h06D:  rddata <= 12'd175;
        9'h06E:  rddata <= 12'd172;
        9'h06F:  rddata <= 12'd169;
        9'h070:  rddata <= 12'd167;
        9'h071:  rddata <= 12'd164;
        9'h072:  rddata <= 12'd161;
        9'h073:  rddata <= 12'd159;
        9'h074:  rddata <= 12'd156;
        9'h075:  rddata <= 12'd153;
        9'h076:  rddata <= 12'd151;
        9'h077:  rddata <= 12'd148;
        9'h078:  rddata <= 12'd146;
        9'h079:  rddata <= 12'd143;
        9'h07A:  rddata <= 12'd141;
        9'h07B:  rddata <= 12'd138;
        9'h07C:  rddata <= 12'd136;
        9'h07D:  rddata <= 12'd134;
        9'h07E:  rddata <= 12'd131;
        9'h07F:  rddata <= 12'd129;
        9'h080:  rddata <= 12'd127;
        9'h081:  rddata <= 12'd125;
        9'h082:  rddata <= 12'd122;
        9'h083:  rddata <= 12'd120;
        9'h084:  rddata <= 12'd118;
        9'h085:  rddata <= 12'd116;
        9'h086:  rddata <= 12'd114;
        9'h087:  rddata <= 12'd112;
        9'h088:  rddata <= 12'd110;
        9'h089:  rddata <= 12'd108;
        9'h08A:  rddata <= 12'd106;
        9'h08B:  rddata <= 12'd104;
        9'h08C:  rddata <= 12'd102;
        9'h08D:  rddata <= 12'd100;
        9'h08E:  rddata <= 12'd98;
        9'h08F:  rddata <= 12'd96;
        9'h090:  rddata <= 12'd94;
        9'h091:  rddata <= 12'd92;
        9'h092:  rddata <= 12'd91;
        9'h093:  rddata <= 12'd89;
        9'h094:  rddata <= 12'd87;
        9'h095:  rddata <= 12'd85;
        9'h096:  rddata <= 12'd83;
        9'h097:  rddata <= 12'd82;
        9'h098:  rddata <= 12'd80;
        9'h099:  rddata <= 12'd78;
        9'h09A:  rddata <= 12'd77;
        9'h09B:  rddata <= 12'd75;
        9'h09C:  rddata <= 12'd74;
        9'h09D:  rddata <= 12'd72;
        9'h09E:  rddata <= 12'd70;
        9'h09F:  rddata <= 12'd69;
        9'h0A0:  rddata <= 12'd67;
        9'h0A1:  rddata <= 12'd66;
        9'h0A2:  rddata <= 12'd64;
        9'h0A3:  rddata <= 12'd63;
        9'h0A4:  rddata <= 12'd62;
        9'h0A5:  rddata <= 12'd60;
        9'h0A6:  rddata <= 12'd59;
        9'h0A7:  rddata <= 12'd57;
        9'h0A8:  rddata <= 12'd56;
        9'h0A9:  rddata <= 12'd55;
        9'h0AA:  rddata <= 12'd53;
        9'h0AB:  rddata <= 12'd52;
        9'h0AC:  rddata <= 12'd51;
        9'h0AD:  rddata <= 12'd49;
        9'h0AE:  rddata <= 12'd48;
        9'h0AF:  rddata <= 12'd47;
        9'h0B0:  rddata <= 12'd46;
        9'h0B1:  rddata <= 12'd45;
        9'h0B2:  rddata <= 12'd43;
        9'h0B3:  rddata <= 12'd42;
        9'h0B4:  rddata <= 12'd41;
        9'h0B5:  rddata <= 12'd40;
        9'h0B6:  rddata <= 12'd39;
        9'h0B7:  rddata <= 12'd38;
        9'h0B8:  rddata <= 12'd37;
        9'h0B9:  rddata <= 12'd36;
        9'h0BA:  rddata <= 12'd35;
        9'h0BB:  rddata <= 12'd34;
        9'h0BC:  rddata <= 12'd33;
        9'h0BD:  rddata <= 12'd32;
        9'h0BE:  rddata <= 12'd31;
        9'h0BF:  rddata <= 12'd30;
        9'h0C0:  rddata <= 12'd29;
        9'h0C1:  rddata <= 12'd28;
        9'h0C2:  rddata <= 12'd27;
        9'h0C3:  rddata <= 12'd26;
        9'h0C4:  rddata <= 12'd25;
        9'h0C5:  rddata <= 12'd24;
        9'h0C6:  rddata <= 12'd23;
        9'h0C7:  rddata <= 12'd23;
        9'h0C8:  rddata <= 12'd22;
        9'h0C9:  rddata <= 12'd21;
        9'h0CA:  rddata <= 12'd20;
        9'h0CB:  rddata <= 12'd20;
        9'h0CC:  rddata <= 12'd19;
        9'h0CD:  rddata <= 12'd18;
        9'h0CE:  rddata <= 12'd17;
        9'h0CF:  rddata <= 12'd17;
        9'h0D0:  rddata <= 12'd16;
        9'h0D1:  rddata <= 12'd15;
        9'h0D2:  rddata <= 12'd15;
        9'h0D3:  rddata <= 12'd14;
        9'h0D4:  rddata <= 12'd13;
        9'h0D5:  rddata <= 12'd13;
        9'h0D6:  rddata <= 12'd12;
        9'h0D7:  rddata <= 12'd12;
        9'h0D8:  rddata <= 12'd11;
        9'h0D9:  rddata <= 12'd10;
        9'h0DA:  rddata <= 12'd10;
        9'h0DB:  rddata <= 12'd9;
        9'h0DC:  rddata <= 12'd9;
        9'h0DD:  rddata <= 12'd8;
        9'h0DE:  rddata <= 12'd8;
        9'h0DF:  rddata <= 12'd7;
        9'h0E0:  rddata <= 12'd7;
        9'h0E1:  rddata <= 12'd7;
        9'h0E2:  rddata <= 12'd6;
        9'h0E3:  rddata <= 12'd6;
        9'h0E4:  rddata <= 12'd5;
        9'h0E5:  rddata <= 12'd5;
        9'h0E6:  rddata <= 12'd5;
        9'h0E7:  rddata <= 12'd4;
        9'h0E8:  rddata <= 12'd4;
        9'h0E9:  rddata <= 12'd4;
        9'h0EA:  rddata <= 12'd3;
        9'h0EB:  rddata <= 12'd3;
        9'h0EC:  rddata <= 12'd3;
        9'h0ED:  rddata <= 12'd2;
        9'h0EE:  rddata <= 12'd2;
        9'h0EF:  rddata <= 12'd2;
        9'h0F0:  rddata <= 12'd2;
        9'h0F1:  rddata <= 12'd1;
        9'h0F2:  rddata <= 12'd1;
        9'h0F3:  rddata <= 12'd1;
        9'h0F4:  rddata <= 12'd1;
        9'h0F5:  rddata <= 12'd1;
        9'h0F6:  rddata <= 12'd1;
        9'h0F7:  rddata <= 12'd1;
        9'h0F8:  rddata <= 12'd0;
        9'h0F9:  rddata <= 12'd0;
        9'h0FA:  rddata <= 12'd0;
        9'h0FB:  rddata <= 12'd0;
        9'h0FC:  rddata <= 12'd0;
        9'h0FD:  rddata <= 12'd0;
        9'h0FE:  rddata <= 12'd0;
        9'h0FF:  rddata <= 12'd0;
        9'h100:  rddata <= 12'd0;
        9'h101:  rddata <= 12'd3;
        9'h102:  rddata <= 12'd6;
        9'h103:  rddata <= 12'd8;
        9'h104:  rddata <= 12'd11;
        9'h105:  rddata <= 12'd14;
        9'h106:  rddata <= 12'd17;
        9'h107:  rddata <= 12'd20;
        9'h108:  rddata <= 12'd22;
        9'h109:  rddata <= 12'd25;
        9'h10A:  rddata <= 12'd28;
        9'h10B:  rddata <= 12'd31;
        9'h10C:  rddata <= 12'd34;
        9'h10D:  rddata <= 12'd37;
        9'h10E:  rddata <= 12'd40;
        9'h10F:  rddata <= 12'd42;
        9'h110:  rddata <= 12'd45;
        9'h111:  rddata <= 12'd48;
        9'h112:  rddata <= 12'd51;
        9'h113:  rddata <= 12'd54;
        9'h114:  rddata <= 12'd57;
        9'h115:  rddata <= 12'd60;
        9'h116:  rddata <= 12'd63;
        9'h117:  rddata <= 12'd66;
        9'h118:  rddata <= 12'd69;
        9'h119:  rddata <= 12'd72;
        9'h11A:  rddata <= 12'd75;
        9'h11B:  rddata <= 12'd78;
        9'h11C:  rddata <= 12'd81;
        9'h11D:  rddata <= 12'd84;
        9'h11E:  rddata <= 12'd87;
        9'h11F:  rddata <= 12'd90;
        9'h120:  rddata <= 12'd93;
        9'h121:  rddata <= 12'd96;
        9'h122:  rddata <= 12'd99;
        9'h123:  rddata <= 12'd102;
        9'h124:  rddata <= 12'd105;
        9'h125:  rddata <= 12'd108;
        9'h126:  rddata <= 12'd111;
        9'h127:  rddata <= 12'd114;
        9'h128:  rddata <= 12'd117;
        9'h129:  rddata <= 12'd120;
        9'h12A:  rddata <= 12'd123;
        9'h12B:  rddata <= 12'd126;
        9'h12C:  rddata <= 12'd130;
        9'h12D:  rddata <= 12'd133;
        9'h12E:  rddata <= 12'd136;
        9'h12F:  rddata <= 12'd139;
        9'h130:  rddata <= 12'd142;
        9'h131:  rddata <= 12'd145;
        9'h132:  rddata <= 12'd148;
        9'h133:  rddata <= 12'd152;
        9'h134:  rddata <= 12'd155;
        9'h135:  rddata <= 12'd158;
        9'h136:  rddata <= 12'd161;
        9'h137:  rddata <= 12'd164;
        9'h138:  rddata <= 12'd168;
        9'h139:  rddata <= 12'd171;
        9'h13A:  rddata <= 12'd174;
        9'h13B:  rddata <= 12'd177;
        9'h13C:  rddata <= 12'd181;
        9'h13D:  rddata <= 12'd184;
        9'h13E:  rddata <= 12'd187;
        9'h13F:  rddata <= 12'd190;
        9'h140:  rddata <= 12'd194;
        9'h141:  rddata <= 12'd197;
        9'h142:  rddata <= 12'd200;
        9'h143:  rddata <= 12'd204;
        9'h144:  rddata <= 12'd207;
        9'h145:  rddata <= 12'd210;
        9'h146:  rddata <= 12'd214;
        9'h147:  rddata <= 12'd217;
        9'h148:  rddata <= 12'd220;
        9'h149:  rddata <= 12'd224;
        9'h14A:  rddata <= 12'd227;
        9'h14B:  rddata <= 12'd231;
        9'h14C:  rddata <= 12'd234;
        9'h14D:  rddata <= 12'd237;
        9'h14E:  rddata <= 12'd241;
        9'h14F:  rddata <= 12'd244;
        9'h150:  rddata <= 12'd248;
        9'h151:  rddata <= 12'd251;
        9'h152:  rddata <= 12'd255;
        9'h153:  rddata <= 12'd258;
        9'h154:  rddata <= 12'd262;
        9'h155:  rddata <= 12'd265;
        9'h156:  rddata <= 12'd268;
        9'h157:  rddata <= 12'd272;
        9'h158:  rddata <= 12'd276;
        9'h159:  rddata <= 12'd279;
        9'h15A:  rddata <= 12'd283;
        9'h15B:  rddata <= 12'd286;
        9'h15C:  rddata <= 12'd290;
        9'h15D:  rddata <= 12'd293;
        9'h15E:  rddata <= 12'd297;
        9'h15F:  rddata <= 12'd300;
        9'h160:  rddata <= 12'd304;
        9'h161:  rddata <= 12'd308;
        9'h162:  rddata <= 12'd311;
        9'h163:  rddata <= 12'd315;
        9'h164:  rddata <= 12'd318;
        9'h165:  rddata <= 12'd322;
        9'h166:  rddata <= 12'd326;
        9'h167:  rddata <= 12'd329;
        9'h168:  rddata <= 12'd333;
        9'h169:  rddata <= 12'd337;
        9'h16A:  rddata <= 12'd340;
        9'h16B:  rddata <= 12'd344;
        9'h16C:  rddata <= 12'd348;
        9'h16D:  rddata <= 12'd352;
        9'h16E:  rddata <= 12'd355;
        9'h16F:  rddata <= 12'd359;
        9'h170:  rddata <= 12'd363;
        9'h171:  rddata <= 12'd367;
        9'h172:  rddata <= 12'd370;
        9'h173:  rddata <= 12'd374;
        9'h174:  rddata <= 12'd378;
        9'h175:  rddata <= 12'd382;
        9'h176:  rddata <= 12'd385;
        9'h177:  rddata <= 12'd389;
        9'h178:  rddata <= 12'd393;
        9'h179:  rddata <= 12'd397;
        9'h17A:  rddata <= 12'd401;
        9'h17B:  rddata <= 12'd405;
        9'h17C:  rddata <= 12'd409;
        9'h17D:  rddata <= 12'd412;
        9'h17E:  rddata <= 12'd416;
        9'h17F:  rddata <= 12'd420;
        9'h180:  rddata <= 12'd424;
        9'h181:  rddata <= 12'd428;
        9'h182:  rddata <= 12'd432;
        9'h183:  rddata <= 12'd436;
        9'h184:  rddata <= 12'd440;
        9'h185:  rddata <= 12'd444;
        9'h186:  rddata <= 12'd448;
        9'h187:  rddata <= 12'd452;
        9'h188:  rddata <= 12'd456;
        9'h189:  rddata <= 12'd460;
        9'h18A:  rddata <= 12'd464;
        9'h18B:  rddata <= 12'd468;
        9'h18C:  rddata <= 12'd472;
        9'h18D:  rddata <= 12'd476;
        9'h18E:  rddata <= 12'd480;
        9'h18F:  rddata <= 12'd484;
        9'h190:  rddata <= 12'd488;
        9'h191:  rddata <= 12'd492;
        9'h192:  rddata <= 12'd496;
        9'h193:  rddata <= 12'd501;
        9'h194:  rddata <= 12'd505;
        9'h195:  rddata <= 12'd509;
        9'h196:  rddata <= 12'd513;
        9'h197:  rddata <= 12'd517;
        9'h198:  rddata <= 12'd521;
        9'h199:  rddata <= 12'd526;
        9'h19A:  rddata <= 12'd530;
        9'h19B:  rddata <= 12'd534;
        9'h19C:  rddata <= 12'd538;
        9'h19D:  rddata <= 12'd542;
        9'h19E:  rddata <= 12'd547;
        9'h19F:  rddata <= 12'd551;
        9'h1A0:  rddata <= 12'd555;
        9'h1A1:  rddata <= 12'd560;
        9'h1A2:  rddata <= 12'd564;
        9'h1A3:  rddata <= 12'd568;
        9'h1A4:  rddata <= 12'd572;
        9'h1A5:  rddata <= 12'd577;
        9'h1A6:  rddata <= 12'd581;
        9'h1A7:  rddata <= 12'd585;
        9'h1A8:  rddata <= 12'd590;
        9'h1A9:  rddata <= 12'd594;
        9'h1AA:  rddata <= 12'd599;
        9'h1AB:  rddata <= 12'd603;
        9'h1AC:  rddata <= 12'd607;
        9'h1AD:  rddata <= 12'd612;
        9'h1AE:  rddata <= 12'd616;
        9'h1AF:  rddata <= 12'd621;
        9'h1B0:  rddata <= 12'd625;
        9'h1B1:  rddata <= 12'd630;
        9'h1B2:  rddata <= 12'd634;
        9'h1B3:  rddata <= 12'd639;
        9'h1B4:  rddata <= 12'd643;
        9'h1B5:  rddata <= 12'd648;
        9'h1B6:  rddata <= 12'd652;
        9'h1B7:  rddata <= 12'd657;
        9'h1B8:  rddata <= 12'd661;
        9'h1B9:  rddata <= 12'd666;
        9'h1BA:  rddata <= 12'd670;
        9'h1BB:  rddata <= 12'd675;
        9'h1BC:  rddata <= 12'd680;
        9'h1BD:  rddata <= 12'd684;
        9'h1BE:  rddata <= 12'd689;
        9'h1BF:  rddata <= 12'd693;
        9'h1C0:  rddata <= 12'd698;
        9'h1C1:  rddata <= 12'd703;
        9'h1C2:  rddata <= 12'd708;
        9'h1C3:  rddata <= 12'd712;
        9'h1C4:  rddata <= 12'd717;
        9'h1C5:  rddata <= 12'd722;
        9'h1C6:  rddata <= 12'd726;
        9'h1C7:  rddata <= 12'd731;
        9'h1C8:  rddata <= 12'd736;
        9'h1C9:  rddata <= 12'd741;
        9'h1CA:  rddata <= 12'd745;
        9'h1CB:  rddata <= 12'd750;
        9'h1CC:  rddata <= 12'd755;
        9'h1CD:  rddata <= 12'd760;
        9'h1CE:  rddata <= 12'd765;
        9'h1CF:  rddata <= 12'd770;
        9'h1D0:  rddata <= 12'd774;
        9'h1D1:  rddata <= 12'd779;
        9'h1D2:  rddata <= 12'd784;
        9'h1D3:  rddata <= 12'd789;
        9'h1D4:  rddata <= 12'd794;
        9'h1D5:  rddata <= 12'd799;
        9'h1D6:  rddata <= 12'd804;
        9'h1D7:  rddata <= 12'd809;
        9'h1D8:  rddata <= 12'd814;
        9'h1D9:  rddata <= 12'd819;
        9'h1DA:  rddata <= 12'd824;
        9'h1DB:  rddata <= 12'd829;
        9'h1DC:  rddata <= 12'd834;
        9'h1DD:  rddata <= 12'd839;
        9'h1DE:  rddata <= 12'd844;
        9'h1DF:  rddata <= 12'd849;
        9'h1E0:  rddata <= 12'd854;
        9'h1E1:  rddata <= 12'd859;
        9'h1E2:  rddata <= 12'd864;
        9'h1E3:  rddata <= 12'd869;
        9'h1E4:  rddata <= 12'd874;
        9'h1E5:  rddata <= 12'd880;
        9'h1E6:  rddata <= 12'd885;
        9'h1E7:  rddata <= 12'd890;
        9'h1E8:  rddata <= 12'd895;
        9'h1E9:  rddata <= 12'd900;
        9'h1EA:  rddata <= 12'd906;
        9'h1EB:  rddata <= 12'd911;
        9'h1EC:  rddata <= 12'd916;
        9'h1ED:  rddata <= 12'd921;
        9'h1EE:  rddata <= 12'd927;
        9'h1EF:  rddata <= 12'd932;
        9'h1F0:  rddata <= 12'd937;
        9'h1F1:  rddata <= 12'd942;
        9'h1F2:  rddata <= 12'd948;
        9'h1F3:  rddata <= 12'd953;
        9'h1F4:  rddata <= 12'd959;
        9'h1F5:  rddata <= 12'd964;
        9'h1F6:  rddata <= 12'd969;
        9'h1F7:  rddata <= 12'd975;
        9'h1F8:  rddata <= 12'd980;
        9'h1F9:  rddata <= 12'd986;
        9'h1FA:  rddata <= 12'd991;
        9'h1FB:  rddata <= 12'd996;
        9'h1FC:  rddata <= 12'd1002;
        9'h1FD:  rddata <= 12'd1007;
        9'h1FE:  rddata <= 12'd1013;
        9'h1FF:  rddata <= 12'd1018;
        default: rddata <= 12'd0;
    endcase

endmodule
