`default_nettype none
`timescale 1 ns / 1 ps

(* rom_style = "distributed" *)
module lut_exp(
    input  wire        clk,
    input  wire  [7:0] addr,
    output reg   [9:0] rddata
);

    always @(posedge clk) case (addr)
        8'h00: rddata <= 10'd0;
        8'h01: rddata <= 10'd3;
        8'h02: rddata <= 10'd6;
        8'h03: rddata <= 10'd8;
        8'h04: rddata <= 10'd11;
        8'h05: rddata <= 10'd14;
        8'h06: rddata <= 10'd17;
        8'h07: rddata <= 10'd20;
        8'h08: rddata <= 10'd22;
        8'h09: rddata <= 10'd25;
        8'h0A: rddata <= 10'd28;
        8'h0B: rddata <= 10'd31;
        8'h0C: rddata <= 10'd34;
        8'h0D: rddata <= 10'd37;
        8'h0E: rddata <= 10'd40;
        8'h0F: rddata <= 10'd42;
        8'h10: rddata <= 10'd45;
        8'h11: rddata <= 10'd48;
        8'h12: rddata <= 10'd51;
        8'h13: rddata <= 10'd54;
        8'h14: rddata <= 10'd57;
        8'h15: rddata <= 10'd60;
        8'h16: rddata <= 10'd63;
        8'h17: rddata <= 10'd66;
        8'h18: rddata <= 10'd69;
        8'h19: rddata <= 10'd72;
        8'h1A: rddata <= 10'd75;
        8'h1B: rddata <= 10'd78;
        8'h1C: rddata <= 10'd81;
        8'h1D: rddata <= 10'd84;
        8'h1E: rddata <= 10'd87;
        8'h1F: rddata <= 10'd90;
        8'h20: rddata <= 10'd93;
        8'h21: rddata <= 10'd96;
        8'h22: rddata <= 10'd99;
        8'h23: rddata <= 10'd102;
        8'h24: rddata <= 10'd105;
        8'h25: rddata <= 10'd108;
        8'h26: rddata <= 10'd111;
        8'h27: rddata <= 10'd114;
        8'h28: rddata <= 10'd117;
        8'h29: rddata <= 10'd120;
        8'h2A: rddata <= 10'd123;
        8'h2B: rddata <= 10'd126;
        8'h2C: rddata <= 10'd130;
        8'h2D: rddata <= 10'd133;
        8'h2E: rddata <= 10'd136;
        8'h2F: rddata <= 10'd139;
        8'h30: rddata <= 10'd142;
        8'h31: rddata <= 10'd145;
        8'h32: rddata <= 10'd148;
        8'h33: rddata <= 10'd152;
        8'h34: rddata <= 10'd155;
        8'h35: rddata <= 10'd158;
        8'h36: rddata <= 10'd161;
        8'h37: rddata <= 10'd164;
        8'h38: rddata <= 10'd168;
        8'h39: rddata <= 10'd171;
        8'h3A: rddata <= 10'd174;
        8'h3B: rddata <= 10'd177;
        8'h3C: rddata <= 10'd181;
        8'h3D: rddata <= 10'd184;
        8'h3E: rddata <= 10'd187;
        8'h3F: rddata <= 10'd190;
        8'h40: rddata <= 10'd194;
        8'h41: rddata <= 10'd197;
        8'h42: rddata <= 10'd200;
        8'h43: rddata <= 10'd204;
        8'h44: rddata <= 10'd207;
        8'h45: rddata <= 10'd210;
        8'h46: rddata <= 10'd214;
        8'h47: rddata <= 10'd217;
        8'h48: rddata <= 10'd220;
        8'h49: rddata <= 10'd224;
        8'h4A: rddata <= 10'd227;
        8'h4B: rddata <= 10'd231;
        8'h4C: rddata <= 10'd234;
        8'h4D: rddata <= 10'd237;
        8'h4E: rddata <= 10'd241;
        8'h4F: rddata <= 10'd244;
        8'h50: rddata <= 10'd248;
        8'h51: rddata <= 10'd251;
        8'h52: rddata <= 10'd255;
        8'h53: rddata <= 10'd258;
        8'h54: rddata <= 10'd262;
        8'h55: rddata <= 10'd265;
        8'h56: rddata <= 10'd268;
        8'h57: rddata <= 10'd272;
        8'h58: rddata <= 10'd276;
        8'h59: rddata <= 10'd279;
        8'h5A: rddata <= 10'd283;
        8'h5B: rddata <= 10'd286;
        8'h5C: rddata <= 10'd290;
        8'h5D: rddata <= 10'd293;
        8'h5E: rddata <= 10'd297;
        8'h5F: rddata <= 10'd300;
        8'h60: rddata <= 10'd304;
        8'h61: rddata <= 10'd308;
        8'h62: rddata <= 10'd311;
        8'h63: rddata <= 10'd315;
        8'h64: rddata <= 10'd318;
        8'h65: rddata <= 10'd322;
        8'h66: rddata <= 10'd326;
        8'h67: rddata <= 10'd329;
        8'h68: rddata <= 10'd333;
        8'h69: rddata <= 10'd337;
        8'h6A: rddata <= 10'd340;
        8'h6B: rddata <= 10'd344;
        8'h6C: rddata <= 10'd348;
        8'h6D: rddata <= 10'd352;
        8'h6E: rddata <= 10'd355;
        8'h6F: rddata <= 10'd359;
        8'h70: rddata <= 10'd363;
        8'h71: rddata <= 10'd367;
        8'h72: rddata <= 10'd370;
        8'h73: rddata <= 10'd374;
        8'h74: rddata <= 10'd378;
        8'h75: rddata <= 10'd382;
        8'h76: rddata <= 10'd385;
        8'h77: rddata <= 10'd389;
        8'h78: rddata <= 10'd393;
        8'h79: rddata <= 10'd397;
        8'h7A: rddata <= 10'd401;
        8'h7B: rddata <= 10'd405;
        8'h7C: rddata <= 10'd409;
        8'h7D: rddata <= 10'd412;
        8'h7E: rddata <= 10'd416;
        8'h7F: rddata <= 10'd420;
        8'h80: rddata <= 10'd424;
        8'h81: rddata <= 10'd428;
        8'h82: rddata <= 10'd432;
        8'h83: rddata <= 10'd436;
        8'h84: rddata <= 10'd440;
        8'h85: rddata <= 10'd444;
        8'h86: rddata <= 10'd448;
        8'h87: rddata <= 10'd452;
        8'h88: rddata <= 10'd456;
        8'h89: rddata <= 10'd460;
        8'h8A: rddata <= 10'd464;
        8'h8B: rddata <= 10'd468;
        8'h8C: rddata <= 10'd472;
        8'h8D: rddata <= 10'd476;
        8'h8E: rddata <= 10'd480;
        8'h8F: rddata <= 10'd484;
        8'h90: rddata <= 10'd488;
        8'h91: rddata <= 10'd492;
        8'h92: rddata <= 10'd496;
        8'h93: rddata <= 10'd501;
        8'h94: rddata <= 10'd505;
        8'h95: rddata <= 10'd509;
        8'h96: rddata <= 10'd513;
        8'h97: rddata <= 10'd517;
        8'h98: rddata <= 10'd521;
        8'h99: rddata <= 10'd526;
        8'h9A: rddata <= 10'd530;
        8'h9B: rddata <= 10'd534;
        8'h9C: rddata <= 10'd538;
        8'h9D: rddata <= 10'd542;
        8'h9E: rddata <= 10'd547;
        8'h9F: rddata <= 10'd551;
        8'hA0: rddata <= 10'd555;
        8'hA1: rddata <= 10'd560;
        8'hA2: rddata <= 10'd564;
        8'hA3: rddata <= 10'd568;
        8'hA4: rddata <= 10'd572;
        8'hA5: rddata <= 10'd577;
        8'hA6: rddata <= 10'd581;
        8'hA7: rddata <= 10'd585;
        8'hA8: rddata <= 10'd590;
        8'hA9: rddata <= 10'd594;
        8'hAA: rddata <= 10'd599;
        8'hAB: rddata <= 10'd603;
        8'hAC: rddata <= 10'd607;
        8'hAD: rddata <= 10'd612;
        8'hAE: rddata <= 10'd616;
        8'hAF: rddata <= 10'd621;
        8'hB0: rddata <= 10'd625;
        8'hB1: rddata <= 10'd630;
        8'hB2: rddata <= 10'd634;
        8'hB3: rddata <= 10'd639;
        8'hB4: rddata <= 10'd643;
        8'hB5: rddata <= 10'd648;
        8'hB6: rddata <= 10'd652;
        8'hB7: rddata <= 10'd657;
        8'hB8: rddata <= 10'd661;
        8'hB9: rddata <= 10'd666;
        8'hBA: rddata <= 10'd670;
        8'hBB: rddata <= 10'd675;
        8'hBC: rddata <= 10'd680;
        8'hBD: rddata <= 10'd684;
        8'hBE: rddata <= 10'd689;
        8'hBF: rddata <= 10'd693;
        8'hC0: rddata <= 10'd698;
        8'hC1: rddata <= 10'd703;
        8'hC2: rddata <= 10'd708;
        8'hC3: rddata <= 10'd712;
        8'hC4: rddata <= 10'd717;
        8'hC5: rddata <= 10'd722;
        8'hC6: rddata <= 10'd726;
        8'hC7: rddata <= 10'd731;
        8'hC8: rddata <= 10'd736;
        8'hC9: rddata <= 10'd741;
        8'hCA: rddata <= 10'd745;
        8'hCB: rddata <= 10'd750;
        8'hCC: rddata <= 10'd755;
        8'hCD: rddata <= 10'd760;
        8'hCE: rddata <= 10'd765;
        8'hCF: rddata <= 10'd770;
        8'hD0: rddata <= 10'd774;
        8'hD1: rddata <= 10'd779;
        8'hD2: rddata <= 10'd784;
        8'hD3: rddata <= 10'd789;
        8'hD4: rddata <= 10'd794;
        8'hD5: rddata <= 10'd799;
        8'hD6: rddata <= 10'd804;
        8'hD7: rddata <= 10'd809;
        8'hD8: rddata <= 10'd814;
        8'hD9: rddata <= 10'd819;
        8'hDA: rddata <= 10'd824;
        8'hDB: rddata <= 10'd829;
        8'hDC: rddata <= 10'd834;
        8'hDD: rddata <= 10'd839;
        8'hDE: rddata <= 10'd844;
        8'hDF: rddata <= 10'd849;
        8'hE0: rddata <= 10'd854;
        8'hE1: rddata <= 10'd859;
        8'hE2: rddata <= 10'd864;
        8'hE3: rddata <= 10'd869;
        8'hE4: rddata <= 10'd874;
        8'hE5: rddata <= 10'd880;
        8'hE6: rddata <= 10'd885;
        8'hE7: rddata <= 10'd890;
        8'hE8: rddata <= 10'd895;
        8'hE9: rddata <= 10'd900;
        8'hEA: rddata <= 10'd906;
        8'hEB: rddata <= 10'd911;
        8'hEC: rddata <= 10'd916;
        8'hED: rddata <= 10'd921;
        8'hEE: rddata <= 10'd927;
        8'hEF: rddata <= 10'd932;
        8'hF0: rddata <= 10'd937;
        8'hF1: rddata <= 10'd942;
        8'hF2: rddata <= 10'd948;
        8'hF3: rddata <= 10'd953;
        8'hF4: rddata <= 10'd959;
        8'hF5: rddata <= 10'd964;
        8'hF6: rddata <= 10'd969;
        8'hF7: rddata <= 10'd975;
        8'hF8: rddata <= 10'd980;
        8'hF9: rddata <= 10'd986;
        8'hFA: rddata <= 10'd991;
        8'hFB: rddata <= 10'd996;
        8'hFC: rddata <= 10'd1002;
        8'hFD: rddata <= 10'd1007;
        8'hFE: rddata <= 10'd1013;
        8'hFF: rddata <= 10'd1018;
        default: rddata <= 10'd0;
    endcase

endmodule
